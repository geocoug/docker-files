netcdf edu_calpoly_marine_morro_bay_met {
dimensions:
	time = 40970 ;
variables:
	int crs ;
		crs:_Storage = "contiguous" ;
		crs:_Endianness = "little" ;
	double time(time) ;
		time:units = "seconds since 1970-01-01T00:00:00Z" ;
		time:standard_name = "time" ;
		time:axis = "T" ;
		time:_ChunkSizes = 40794 ;
		time:_CoordinateAxisType = "Time" ;
		time:actual_range = 1454284800., 1571962037. ;
		time:calendar = "gregorian" ;
		time:ioos_category = "Time" ;
		time:long_name = "Time" ;
		time:time_origin = "01-JAN-1970 00:00:00" ;
		time:_Storage = "contiguous" ;
		time:_Endianness = "little" ;
	string station ;
		station:cf_role = "timeseries_id" ;
		station:long_name = "Morro Bay - BS1 MET" ;
		station:_Encoding = "ISO-8859-1" ;
		station:ioos_category = "Identifier" ;
		station:ioos_code = "urn:ioos:station:com.axiomdatascience:57163" ;
		station:short_name = "edu_calpoly_marine_morro_bay_met" ;
		station:type = "fixed" ;
		station:_Storage = "contiguous" ;
	double latitude ;
		latitude:axis = "Y" ;
		latitude:_CoordinateAxisType = "Lat" ;
		latitude:actual_range = 35.33382, 35.33382 ;
		latitude:ioos_category = "Location" ;
		latitude:long_name = "Latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:_Storage = "contiguous" ;
		latitude:_Endianness = "little" ;
	double longitude ;
		longitude:axis = "X" ;
		longitude:_CoordinateAxisType = "Lon" ;
		longitude:actual_range = -120.84725, -120.84725 ;
		longitude:ioos_category = "Location" ;
		longitude:long_name = "Longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:_Storage = "contiguous" ;
		longitude:_Endianness = "little" ;
	double z ;
		z:_FillValue = -9999.9 ;
		z:axis = "Z" ;
		z:_ChunkSizes = 1 ;
		z:_CoordinateAxisType = "Height" ;
		z:_CoordinateZisPositive = "up" ;
		z:actual_range = 0., 0. ;
		z:ioos_category = "Location" ;
		z:least_significant_digit = 2. ;
		z:long_name = "Altitude" ;
		z:positive = "up" ;
		z:standard_name = "altitude" ;
		z:units = "m" ;
		z:_Storage = "contiguous" ;
		z:_Endianness = "little" ;
	double air_temperature(time) ;
		air_temperature:_FillValue = -9999.9 ;
		air_temperature:_ChunkSizes = 40794, 1 ;
		air_temperature:actual_range = -9.35, 34.03 ;
		air_temperature:id = "1000293" ;
		air_temperature:ioos_category = "Other" ;
		air_temperature:long_name = "Air Temperature" ;
		air_temperature:platform = "station" ;
		air_temperature:standard_name = "air_temperature" ;
		air_temperature:standard_name_url = "http://mmisw.org/ont/cf/parameter/air_temperature" ;
		air_temperature:units = "degree_Celsius" ;
		air_temperature:coordinates = "time z longitude latitude" ;
		air_temperature:_Storage = "chunked" ;
		air_temperature:_ChunkSizes = 40970 ;
		air_temperature:_Shuffle = "true" ;
		air_temperature:_DeflateLevel = 1 ;
		air_temperature:_Endianness = "little" ;
	double air_pressure(time) ;
		air_pressure:_FillValue = -9999.9 ;
		air_pressure:_ChunkSizes = 40794, 1 ;
		air_pressure:actual_range = 990.38, 1031.56 ;
		air_pressure:id = "1000289" ;
		air_pressure:ioos_category = "Other" ;
		air_pressure:long_name = "Barometric Pressure" ;
		air_pressure:platform = "station" ;
		air_pressure:standard_name = "air_pressure" ;
		air_pressure:standard_name_url = "http://mmisw.org/ont/cf/parameter/air_pressure" ;
		air_pressure:units = "millibars" ;
		air_pressure:coordinates = "time z longitude latitude" ;
		air_pressure:_Storage = "chunked" ;
		air_pressure:_ChunkSizes = 40970 ;
		air_pressure:_Shuffle = "true" ;
		air_pressure:_DeflateLevel = 1 ;
		air_pressure:_Endianness = "little" ;
	double dew_point_temperature(time) ;
		dew_point_temperature:_FillValue = -9999.9 ;
		dew_point_temperature:_ChunkSizes = 40794, 1 ;
		dew_point_temperature:actual_range = -19.15, 34.03 ;
		dew_point_temperature:id = "1000290" ;
		dew_point_temperature:ioos_category = "Other" ;
		dew_point_temperature:long_name = "Dew Point" ;
		dew_point_temperature:platform = "station" ;
		dew_point_temperature:standard_name = "dew_point_temperature" ;
		dew_point_temperature:standard_name_url = "http://mmisw.org/ont/cf/parameter/dew_point_temperature" ;
		dew_point_temperature:units = "degree_Celsius" ;
		dew_point_temperature:coordinates = "time z longitude latitude" ;
		dew_point_temperature:_Storage = "chunked" ;
		dew_point_temperature:_ChunkSizes = 40970 ;
		dew_point_temperature:_Shuffle = "true" ;
		dew_point_temperature:_DeflateLevel = 1 ;
		dew_point_temperature:_Endianness = "little" ;
	double lwe_precipitation_rate_cm_time__sum_over_pt2m(time) ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:_FillValue = -9999.9 ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:_ChunkSizes = 40794, 1 ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:actual_range = 0., 21.5 ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:cell_methods = "time: sum" ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:id = "1000215" ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:interval = "PT2M" ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:ioos_category = "Other" ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:long_name = "Precipitation (increment)" ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:platform = "station" ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:standard_name = "lwe_precipitation_rate" ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:standard_name_url = "http://mmisw.org/ont/cf/parameter/lwe_precipitation_rate" ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:units = "mm" ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:coordinates = "time z longitude latitude" ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:_Storage = "chunked" ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:_ChunkSizes = 40970 ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:_Shuffle = "true" ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:_DeflateLevel = 1 ;
		lwe_precipitation_rate_cm_time__sum_over_pt2m:_Endianness = "little" ;
	double relative_humidity(time) ;
		relative_humidity:_FillValue = -9999.9 ;
		relative_humidity:_ChunkSizes = 40794, 1 ;
		relative_humidity:actual_range = 0., 100. ;
		relative_humidity:id = "1000291" ;
		relative_humidity:ioos_category = "Other" ;
		relative_humidity:long_name = "Relative Humidity" ;
		relative_humidity:platform = "station" ;
		relative_humidity:standard_name = "relative_humidity" ;
		relative_humidity:standard_name_url = "http://mmisw.org/ont/cf/parameter/relative_humidity" ;
		relative_humidity:units = "%" ;
		relative_humidity:coordinates = "time z longitude latitude" ;
		relative_humidity:_Storage = "chunked" ;
		relative_humidity:_ChunkSizes = 40970 ;
		relative_humidity:_Shuffle = "true" ;
		relative_humidity:_DeflateLevel = 1 ;
		relative_humidity:_Endianness = "little" ;
	double solar_irradiance(time) ;
		solar_irradiance:_FillValue = -9999.9 ;
		solar_irradiance:_ChunkSizes = 40794, 1 ;
		solar_irradiance:actual_range = 0., 892.81 ;
		solar_irradiance:id = "1000292" ;
		solar_irradiance:ioos_category = "Other" ;
		solar_irradiance:long_name = "Solar Radiation" ;
		solar_irradiance:platform = "station" ;
		solar_irradiance:standard_name = "solar_irradiance" ;
		solar_irradiance:standard_name_url = "http://mmisw.org/ont/cf/parameter/solar_irradiance" ;
		solar_irradiance:units = "W.m-2" ;
		solar_irradiance:coordinates = "time z longitude latitude" ;
		solar_irradiance:_Storage = "chunked" ;
		solar_irradiance:_ChunkSizes = 40970 ;
		solar_irradiance:_Shuffle = "true" ;
		solar_irradiance:_DeflateLevel = 1 ;
		solar_irradiance:_Endianness = "little" ;
	double wind_chill_temperature(time) ;
		wind_chill_temperature:_FillValue = -9999.9 ;
		wind_chill_temperature:_ChunkSizes = 40794, 1 ;
		wind_chill_temperature:actual_range = -19.15, 34.03 ;
		wind_chill_temperature:id = "1000294" ;
		wind_chill_temperature:ioos_category = "Other" ;
		wind_chill_temperature:long_name = "Wind Chill" ;
		wind_chill_temperature:platform = "station" ;
		wind_chill_temperature:standard_name = "wind_chill_temperature" ;
		wind_chill_temperature:standard_name_url = "http://mmisw.org/ont/unknown/parameter/wind_chill_temperature" ;
		wind_chill_temperature:units = "degree_Celsius" ;
		wind_chill_temperature:coordinates = "time z longitude latitude" ;
		wind_chill_temperature:_Storage = "chunked" ;
		wind_chill_temperature:_ChunkSizes = 40970 ;
		wind_chill_temperature:_Shuffle = "true" ;
		wind_chill_temperature:_DeflateLevel = 1 ;
		wind_chill_temperature:_Endianness = "little" ;
	double wind_speed(time) ;
		wind_speed:_FillValue = -9999.9 ;
		wind_speed:_ChunkSizes = 40794, 1 ;
		wind_speed:actual_range = 0., 18.01 ;
		wind_speed:id = "1000296" ;
		wind_speed:ioos_category = "Other" ;
		wind_speed:long_name = "Wind Speed" ;
		wind_speed:platform = "station" ;
		wind_speed:standard_name = "wind_speed" ;
		wind_speed:standard_name_url = "http://mmisw.org/ont/cf/parameter/wind_speed" ;
		wind_speed:units = "m.s-1" ;
		wind_speed:coordinates = "time z longitude latitude" ;
		wind_speed:_Storage = "chunked" ;
		wind_speed:_ChunkSizes = 40970 ;
		wind_speed:_Shuffle = "true" ;
		wind_speed:_DeflateLevel = 1 ;
		wind_speed:_Endianness = "little" ;
	double wind_from_direction(time) ;
		wind_from_direction:_FillValue = -9999.9 ;
		wind_from_direction:_ChunkSizes = 40794, 1 ;
		wind_from_direction:actual_range = 0.04, 359.88 ;
		wind_from_direction:id = "1000295" ;
		wind_from_direction:ioos_category = "Other" ;
		wind_from_direction:long_name = "Wind From Direction" ;
		wind_from_direction:platform = "station" ;
		wind_from_direction:standard_name = "wind_from_direction" ;
		wind_from_direction:standard_name_url = "http://mmisw.org/ont/cf/parameter/wind_from_direction" ;
		wind_from_direction:units = "degrees" ;
		wind_from_direction:coordinates = "time z longitude latitude" ;
		wind_from_direction:_Storage = "chunked" ;
		wind_from_direction:_ChunkSizes = 40970 ;
		wind_from_direction:_Shuffle = "true" ;
		wind_from_direction:_DeflateLevel = 1 ;
		wind_from_direction:_Endianness = "little" ;

// global attributes:
		:Conventions = "IOOS-1.2, CF-1.6, ACDD-1.3" ;
		:date_created = "2020-04-22T22:29:00Z" ;
		:featureType = "TimeSeries" ;
		:cdm_data_type = "TimeSeries" ;
		:acknowledgment = "Data collection was supported by multiple awards to California Polytechnic State University and an award from NOAA\'s Integrated Observing System to the Central and Northern California Ocean Observing System at the Monterey Bay Aquarium Research Institute (NA11NOS0120032)." ;
		:cdm_timeseries_variables = "station,longitude,latitude" ;
		:comment = "Data produced by Ryan Walter with partial funding from CeNCOOS (cencoos_communicatons@mbari.org)" ;
		:contributor_email = "cencoos_communications@mbari.org,feedback@axiomdatascience.com" ;
		:contributor_name = "Central & Northern California Ocean Observing System (CeNCOOS),Axiom Data Science" ;
		:contributor_role = "contributor,processor" ;
		:contributor_role_vocabulary = "NERC" ;
		:contributor_url = "http://cencoos.org/,https://www.axiomdatascience.com" ;
		:coverage_content_type = "physicalMeasurement" ;
		:creator_country = "USA" ;
		:creator_email = "rkwalter@calpoly.edu" ;
		:creator_institution = "California Polytechnic State University, San Luis Obispo" ;
		:creator_name = "Ryan Walter" ;
		:creator_role = "pi" ;
		:creator_sector = "academic" ;
		:creator_type = "person" ;
		:creator_url = "http://www.marine.calpoly.edu" ;
		:Easternmost_Easting = -120.84725 ;
		:geospatial_lat_max = 35.33382 ;
		:geospatial_lat_min = 35.33382 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_max = -120.84725 ;
		:geospatial_lon_min = -120.84725 ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_vertical_positive = "up" ;
		:geospatial_vertical_units = "m" ;
		:history = "Downloaded from California Polytechnic State University, Center for Coastal Marine Sciences at http://cpool1.marine.calpoly.edu/cpool/CCMS_MorroBay/\n2020-04-22T22:22:19Z http://cpool1.marine.calpoly.edu/cpool/CCMS_MorroBay/\n2020-04-22T22:22:19Z http://erddap.stage.sensors.axds.co/erddap/tabledap/edu_calpoly_marine_morro_bay_met.nc" ;
		:infoUrl = "https://sensors.ioos.us/#metadata/57163/station" ;
		:institution = "California Polytechnic State University, San Luis Obispo" ;
		:instrument = "Nova Lynx 100" ;
		:ISO_Topic_Categories = "Oceans" ;
		:keywords = "Earth Science > Oceans" ;
		:keywords_vocabulary = "GCMD Earth Science Keywords. Version 5.3.3" ;
		:license = "The data may be used and redistributed for free but is not intended\nfor legal use, since it may contain inaccuracies. Neither the data\nContributor, ERD, NOAA, nor the United States Government, nor any\nof their employees or contractors, makes any warranty, express or\nimplied, including warranties of merchantability and fitness for a\nparticular purpose, or assumes any legal liability for the accuracy,\ncompleteness, or usefulness, of this information." ;
		:metadata_conventions = "CF-1.6,ACDD-1.3" ;
		:metadata_link = "http://www.marine.calpoly.edu" ;
		:Northernmost_Northing = 35.33382 ;
		:platform_name = "Morro Bay - BS1 MET" ;
		:platform_vocabulary = "http://mmisw.org/ont/ioos/platform" ;
		:processing_level = "Level 2" ;
		:program = "CeNCOOS" ;
		:project = "CeNCOOS" ;
		:publisher_country = "USA" ;
		:publisher_email = "cencoos_communicatons@mbari.org" ;
		:publisher_institution = "California Polytechnic State University, Center for Coastal Marine Sciences" ;
		:publisher_name = "CeNCOOS" ;
		:publisher_sector = "academic" ;
		:publisher_type = "institution" ;
		:publisher_url = "http://www.cencoos.org" ;
		:references = "http://www.slosea.org/about/dash.php,http://cpool1.marine.calpoly.edu/cpool/CCMS_MorroBay/,https://www.cencoos.org/data/shore/morro," ;
		:sea_name = "NE Pacific" ;
		:source = "Station mounded on a large tripod resting on the sea floor." ;
		:sourceUrl = "http://cpool1.marine.calpoly.edu/cpool/CCMS_MorroBay/" ;
		:Southernmost_Northing = 35.33382 ;
		:standard_name_vocabulary = "CF Standard Name Table v72" ;
		:summary = "Morro Bay BS1 Met station is located in the back of Morro Bay, CA and owned by California Polytechnic State University of San Luis Obispo. The station is mounted on a large tripod, resting on the seafloor. A Nova Lynx 100 Weather Station is fixed at 3 meters above MLLW to a pole extending from the tripod and reports the following in near real-time: wind speed, wind direction, air temperature, barometric pressure, precipitation, relative humidity, and solar radiation. The instrument is maintained and operated by San Luis Obispo Science and Ecosystem Alliance (SLOSEA), a part of the Cal Poly Center for Coastal Marine Sciences." ;
		:time_coverage_end = "2019-10-25T00:07:17Z" ;
		:time_coverage_start = "2016-02-01T00:00:00Z" ;
		:title = "CeNCOOS met monitoring at Morro Bay (BS1)." ;
		:Westernmost_Easting = -120.84725 ;
		:id = "bs1-met" ;
		:naming_authority = "edu.calpoly.marine" ;
		:platform = "morro-bay-bs1-met" ;
		:_NCProperties = "version=2,netcdf=4.6.2,hdf5=1.10.5" ;
		:_SuperblockVersion = 0 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;
data:

 time = 823132800, 823133700, 823134600, 823135500, 823136400, 823137300,
    823138200, 823139100, 823140000, 823140900, 823141800, 823142700,
    823143600, 823144500, 823145400, 823146300, 823147200, 823148100,
    823149000, 823149900, 823150800, 823151700, 823152600, 823153500,
    823154400, 823155300, 823156200, 823157100, 823158000, 823158900,
    823159800, 823160700, 823161600, 823162500, 823163400, 823164300,
    823165200, 823166100, 823167000, 823167900, 823168800, 823169700,
    823170600, 823171500, 823172400, 823173300, 823174200, 823175100,
    823176000, 823176900, 823177800, 823178700, 823179600, 823180500,
    823181400, 823182300, 823183200, 823184100, 823185000, 823185900,
    823186800, 823187700, 823188600, 823189500, 823190400, 823191300,
    823192200, 823193100, 823194000, 823194900, 823195800, 823196700,
    823197600, 823198500, 823199400, 823200300, 823201200, 823202100,
    823203000, 823203900, 823204800, 823205700, 823206600, 823207500,
    823208400, 823209300, 823210200, 823211100, 823212000, 823212900,
    823213800, 823214700, 823215600, 823216500, 823217400, 823218300,
    823219200, 823220100, 823221000, 823221900, 823222800, 823223700,
    823224600, 823225500, 823226400, 823227300, 823228200, 823229100,
    823230000, 823230900, 823231800, 823232700, 823233600, 823234500,
    823235400, 823236300, 823237200, 823238100, 823239000, 823239900,
    823240800, 823241700, 823242600, 823243500, 823244400, 823245300,
    823246200, 823247100, 823248000, 823248900, 823249800, 823250700,
    823251600, 823252500, 823253400, 823254300, 823255200, 823256100,
    823257000, 823257900, 823258800, 823259700, 823260600, 823261500,
    823262400, 823263300, 823264200, 823265100, 823266000, 823266900,
    823267800, 823268700, 823269600, 823270500, 823271400, 823272300,
    823273200, 823274100, 823275000, 823275900, 823276800, 823277700,
    823278600, 823279500, 823280400, 823281300, 823282200, 823283100,
    823284000, 823284900, 823285800, 823286700, 823287600, 823288500,
    823289400, 823290300, 823291200, 823292100, 823293000, 823293900,
    823294800, 823295700, 823296600, 823297500, 823298400, 823299300,
    823300200, 823301100, 823302000, 823302900, 823303800, 823304700,
    823305600, 823306500, 823307400, 823308300, 823309200, 823310100,
    823311000, 823311900, 823312800, 823313700, 823314600, 823315500,
    823316400, 823317300, 823318200, 823319100, 823320000, 823320900,
    823321800, 823322700, 823323600, 823324500, 823325400, 823326300,
    823327200, 823328100, 823329000, 823329900, 823330800, 823331700,
    823332600, 823333500, 823334400, 823335300, 823336200, 823337100,
    823338000, 823338900, 823339800, 823340700, 823341600, 823342500,
    823343400, 823344300, 823345200, 823346100, 823347000, 823347900,
    823348800, 823349700, 823350600, 823351500, 823352400, 823353300,
    823354200, 823355100, 823356000, 823356900, 823357800, 823358700,
    823359600, 823360500, 823361400, 823362300, 823363200, 823364100,
    823365000, 823365900, 823366800, 823367700, 823368600, 823369500,
    823370400, 823371300, 823372200, 823373100, 823374000, 823374900,
    823375800, 823376700, 823377600, 823378500, 823379400, 823380300,
    823381200, 823382100, 823383000, 823383900, 823384800, 823385700,
    823386600, 823387500, 823388400, 823389300, 823390200, 823391100,
    823392000, 823392900, 823393800, 823394700, 823395600, 823396500,
    823397400, 823398300, 823399200, 823400100, 823401000, 823401900,
    823402800, 823403700, 823404600, 823405500, 823406400, 823407300,
    823408200, 823409100, 823410000, 823410900, 823411800, 823412700,
    823413600, 823414500, 823415400, 823416300, 823417200, 823418100,
    823419000, 823419900, 823420800, 823421700, 823422600, 823423500,
    823424400, 823425300, 823426200, 823427100, 823428000, 823428900,
    823429800, 823430700, 823431600, 823432500, 823433400, 823434300,
    823435200, 823436100, 823437000, 823437900, 823438800, 823439700,
    823440600, 823441500, 823442400, 823443300, 823444200, 823445100,
    823446000, 823446900, 823447800, 823448700, 823449600, 823450500,
    823451400, 823452300, 823453200, 823454100, 823455000, 823455900,
    823456800, 823457700, 823458600, 823459500, 823460400, 823461300,
    823462200, 823463100, 823464000, 823464900, 823465800, 823466700,
    823467600, 823468500, 823469400, 823470300, 823471200, 823472100,
    823473000, 823473900, 823474800, 823475700, 823476600, 823477500,
    823478400, 823479300, 823480200, 823481100, 823482000, 823482900,
    823483800, 823484700, 823485600, 823486500, 823487400, 823488300,
    823489200, 823490100, 823491000, 823491900, 823492800, 823493700,
    823494600, 823495500, 823496400, 823497300, 823498200, 823499100,
    823500000, 823500900, 823501800, 823502700, 823503600, 823504500,
    823505400, 823506300, 823507200, 823508100, 823509000, 823509900,
    823510800, 823511700, 823512600, 823513500, 823514400, 823515300,
    823516200, 823517100, 823518000, 823518900, 823519800, 823520700,
    823521600, 823522500, 823523400, 823524300, 823525200, 823526100,
    823527000, 823527900, 823528800, 823529700, 823530600, 823531500,
    823532400, 823533300, 823534200, 823535100, 823536000, 823536900,
    823537800, 823538700, 823539600, 823540500, 823541400, 823542300,
    823543200, 823544100, 823545000, 823545900, 823546800, 823547700,
    823548600, 823549500, 823550400, 823551300, 823552200, 823553100,
    823554000, 823554900, 823555800, 823556700, 823557600, 823558500,
    823559400, 823560300, 823561200, 823562100, 823563000, 823563900,
    823564800, 823565700, 823566600, 823567500, 823568400, 823569300,
    823570200, 823571100, 823572000, 823572900, 823573800, 823574700,
    823575600, 823576500, 823577400, 823578300, 823579200, 823580100,
    823581000, 823581900, 823582800, 823583700, 823584600, 823585500,
    823586400, 823587300, 823588200, 823589100, 823590000, 823590900,
    823591800, 823592700, 823593600, 823594500, 823595400, 823596300,
    823597200, 823598100, 823599000, 823599900, 823600800, 823601700,
    823602600, 823603500, 823604400, 823605300, 823606200, 823607100,
    823608000, 823608900, 823609800, 823610700, 823611600, 823612500,
    823613400, 823614300, 823615200, 823616100, 823617000, 823617900,
    823618800, 823619700, 823620600, 823621500, 823622400, 823623300,
    823624200, 823625100, 823626000, 823626900, 823627800, 823628700,
    823629600, 823630500, 823631400, 823632300, 823633200, 823634100,
    823635000, 823635900, 823636800, 823637700, 823638600, 823639500,
    823640400, 823641300, 823642200, 823643100, 823644000, 823644900,
    823645800, 823646700, 823647600, 823648500, 823649400, 823650300,
    823651200, 823652100, 823653000, 823653900, 823654800, 823655700,
    823656600, 823657500, 823658400, 823659300, 823660200, 823661100,
    823662000, 823662900, 823663800, 823664700, 823665600, 823666500,
    823667400, 823668300, 823669200, 823670100, 823671000, 823671900,
    823672800, 823673700, 823674600, 823675500, 823676400, 823677300,
    823678200, 823679100, 823680000, 823680900, 823681800, 823682700,
    823683600, 823684500, 823685400, 823686300, 823687200, 823688100,
    823689000, 823689900, 823690800, 823691700, 823692600, 823693500,
    823694400, 823695300, 823696200, 823697100, 823698000, 823698900,
    823699800, 823700700, 823701600, 823702500, 823703400, 823704300,
    823705200, 823706100, 823707000, 823707900, 823708800, 823709700,
    823710600, 823711500, 823712400, 823713300, 823714200, 823715100,
    823716000, 823716900, 823717800, 823718700, 823719600, 823720500,
    823721400, 823722300, 823723200, 823724100, 823725000, 823725900,
    823726800, 823727700, 823728600, 823729500, 823730400, 823731300,
    823732200, 823733100, 823734000, 823734900, 823735800, 823736700,
    823737600, 823738500, 823739400, 823740300, 823741200, 823742100,
    823743000, 823743900, 823744800, 823745700, 823746600, 823747500,
    823748400, 823749300, 823750200, 823751100, 823752000, 823752900,
    823753800, 823754700, 823755600, 823756500, 823757400, 823758300,
    823759200, 823760100, 823761000, 823761900, 823762800, 823763700,
    823764600, 823765500, 823766400, 823767300, 823768200, 823769100,
    823770000, 823770900, 823771800, 823772700, 823773600, 823774500,
    823775400, 823776300, 823777200, 823778100, 823779000, 823779900,
    823780800, 823781700, 823782600, 823783500, 823784400, 823785300,
    823786200, 823787100, 823788000, 823788900, 823789800, 823790700,
    823791600, 823792500, 823793400, 823794300, 823795200, 823796100,
    823797000, 823797900, 823798800, 823799700, 823800600, 823801500,
    823802400, 823803300, 823804200, 823805100, 823806000, 823806900,
    823807800, 823808700, 823809600, 823810500, 823811400, 823812300,
    823813200, 823814100, 823815000, 823815900, 823816800, 823817700,
    823818600, 823819500, 823820400, 823821300, 823822200, 823823100,
    823824000, 823824900, 823825800, 823826700, 823827600, 823828500,
    823829400, 823830300, 823831200, 823832100, 823833000, 823833900,
    823834800, 823835700, 823836600, 823837500, 823838400, 823839300,
    823840200, 823841100, 823842000, 823842900, 823843800, 823844700,
    823845600, 823846500, 823847400, 823848300, 823849200, 823850100,
    823851000, 823851900, 823852800, 823853700, 823854600, 823855500,
    823856400, 823857300, 823858200, 823859100, 823860000, 823860900,
    823861800, 823862700, 823863600, 823864500, 823865400, 823866300,
    823867200, 823868100, 823869000, 823869900, 823870800, 823871700,
    823872600, 823873500, 823874400, 823875300, 823876200, 823877100,
    823878000, 823878900, 823879800, 823880700, 823881600, 823882500,
    823883400, 823884300, 823885200, 823886100, 823887000, 823887900,
    823888800, 823889700, 823890600, 823891500, 823892400, 823893300,
    823894200, 823895100, 823896000, 823896900, 823897800, 823898700,
    823899600, 823900500, 823901400, 823902300, 823903200, 823904100,
    823905000, 823905900, 823906800, 823907700, 823908600, 823909500,
    823910400, 823911300, 823912200, 823913100, 823914000, 823914900,
    823915800, 823916700, 823917600, 823918500, 823919400, 823920300,
    823921200, 823922100, 823923000, 823923900, 823924800, 823925700,
    823926600, 823927500, 823928400, 823929300, 823930200, 823931100,
    823932000, 823932900, 823933800, 823934700, 823935600, 823936500,
    823937400, 823938300, 823939200, 823940100, 823941000, 823941900,
    823942800, 823943700, 823944600, 823945500, 823946400, 823947300,
    823948200, 823949100, 823950000, 823950900, 823951800, 823952700,
    823953600, 823954500, 823955400, 823956300, 823957200, 823958100,
    823959000, 823959900, 823960800, 823961700, 823962600, 823963500,
    823964400, 823965300, 823966200, 823967100, 823968000, 823968900,
    823969800, 823970700, 823971600, 823972500, 823973400, 823974300,
    823975200, 823976100, 823977000, 823977900, 823978800, 823979700,
    823980600, 823981500, 823982400, 823983300, 823984200, 823985100,
    823986000, 823986900, 823987800, 823988700, 823989600, 823990500,
    823991400, 823992300, 823993200, 823994100, 823995000, 823995900,
    823996800, 823997700, 823998600, 823999500, 824000400, 824001300,
    824002200, 824003100, 824004000, 824004900, 824005800, 824006700,
    824007600, 824008500, 824009400, 824010300, 824011200, 824012100,
    824013000, 824013900, 824014800, 824015700, 824016600, 824017500,
    824018400, 824019300, 824020200, 824021100, 824022000, 824022900,
    824023800, 824024700, 824025600, 824026500, 824027400, 824028300,
    824029200, 824030100, 824031000, 824031900, 824032800, 824033700,
    824034600, 824035500, 824036400, 824037300, 824038200, 824039100,
    824040000, 824040900, 824041800, 824042700, 824043600, 824044500,
    824045400, 824046300, 824047200, 824048100, 824049000, 824049900,
    824050800, 824051700, 824052600, 824053500, 824054400, 824055300,
    824056200, 824057100, 824058000, 824058900, 824059800, 824060700,
    824061600, 824062500, 824063400, 824064300, 824065200, 824066100,
    824067000, 824067900, 824068800, 824069700, 824070600, 824071500,
    824072400, 824073300, 824074200, 824075100, 824076000, 824076900,
    824077800, 824078700, 824079600, 824080500, 824081400, 824082300,
    824083200, 824084100, 824085000, 824085900, 824086800, 824087700,
    824088600, 824089500, 824090400, 824091300, 824092200, 824093100,
    824094000, 824094900, 824095800, 824096700, 824097600, 824098500,
    824099400, 824100300, 824101200, 824102100, 824103000, 824103900,
    824104800, 824105700, 824106600, 824107500, 824108400, 824109300,
    824110200, 824111100, 824112000, 824112900, 824113800, 824114700,
    824115600, 824116500, 824117400, 824118300, 824119200, 824120100,
    824121000, 824121900, 824122800, 824123700, 824124600, 824125500,
    824126400, 824127300, 824128200, 824129100, 824130000, 824130900,
    824131800, 824132700, 824133600, 824134500, 824135400, 824136300,
    824137200, 824138100, 824139000, 824139900, 824140800, 824141700,
    824142600, 824143500, 824144400, 824145300, 824146200, 824147100,
    824148000, 824148900, 824149800, 824150700, 824151600, 824152500,
    824153400, 824154300, 824155200, 824156100, 824157000, 824157900,
    824158800, 824159700, 824160600, 824161500, 824162400, 824163300,
    824164200, 824165100, 824166000, 824166900, 824167800, 824168700,
    824169600, 824170500, 824171400, 824172300, 824173200, 824174100,
    824175000, 824175900, 824176800, 824177700, 824178600, 824179500,
    824180400, 824181300, 824182200, 824183100, 824184000, 824184900,
    824185800, 824186700, 824187600, 824188500, 824189400, 824190300,
    824191200, 824192100, 824193000, 824193900, 824194800, 824195700,
    824196600, 824197500, 824198400, 824199300, 824200200, 824201100,
    824202000, 824202900, 824203800, 824204700, 824205600, 824206500,
    824207400, 824208300, 824209200, 824210100, 824211000, 824211900,
    824212800, 824213700, 824214600, 824215500, 824216400, 824217300,
    824218200, 824219100, 824220000, 824220900, 824221800, 824222700,
    824223600, 824224500, 824225400, 824226300, 824227200, 824228100,
    824229000, 824229900, 824230800, 824231700, 824232600, 824233500,
    824234400, 824235300, 824236200, 824237100, 824238000, 824238900,
    824239800, 824240700, 824241600, 824242500, 824243400, 824244300,
    824245200, 824246100, 824247000, 824247900, 824248800, 824249700,
    824250600, 824251500, 824252400, 824253300, 824254200, 824255100,
    824256000, 824256900, 824257800, 824258700, 824259600, 824260500,
    824261400, 824262300, 824263200, 824264100, 824265000, 824265900,
    824266800, 824267700, 824268600, 824269500, 824270400, 824271300,
    824272200, 824273100, 824274000, 824274900, 824275800, 824276700,
    824277600, 824278500, 824279400, 824280300, 824281200, 824282100,
    824283000, 824283900, 824284800, 824285700, 824286600, 824287500,
    824288400, 824289300, 824290200, 824291100, 824292000, 824292900,
    824293800, 824294700, 824295600, 824296500, 824297400, 824298300,
    824299200, 824300100, 824301000, 824301900, 824302800, 824303700,
    824304600, 824305500, 824306400, 824307300, 824308200, 824309100,
    824310000, 824310900, 824311800, 824312700, 824313600, 824314500,
    824315400, 824316300, 824317200, 824318100, 824319000, 824319900,
    824320800, 824321700, 824322600, 824323500, 824324400, 824325300,
    824326200, 824327100, 824328000, 824328900, 824329800, 824330700,
    824331600, 824332500, 824333400, 824334300, 824335200, 824336100,
    824337000, 824337900, 824338800, 824339700, 824340600, 824341500,
    824342400, 824343300, 824344200, 824345100, 824346000, 824346900,
    824347800, 824348700, 824349600, 824350500, 824351400, 824352300,
    824353200, 824354100, 824355000, 824355900, 824356800, 824357700,
    824358600, 824359500, 824360400, 824361300, 824362200, 824363100,
    824364000, 824364900, 824365800, 824366700, 824367600, 824368500,
    824369400, 824370300, 824371200, 824372100, 824373000, 824373900,
    824374800, 824375700, 824376600, 824377500, 824378400, 824379300,
    824380200, 824381100, 824382000, 824382900, 824383800, 824384700,
    824385600, 824386500, 824387400, 824388300, 824389200, 824390100,
    824391000, 824391900, 824392800, 824393700, 824394600, 824395500,
    824396400, 824397300, 824398200, 824399100, 824400000, 824400900,
    824401800, 824402700, 824403600, 824404500, 824405400, 824406300,
    824407200, 824408100, 824409000, 824409900, 824410800, 824411700,
    824412600, 824413500, 824414400, 824415300, 824416200, 824417100,
    824418000, 824418900, 824419800, 824420700, 824421600, 824422500,
    824423400, 824424300, 824425200, 824426100, 824427000, 824427900,
    824428800, 824429700, 824430600, 824431500, 824432400, 824433300,
    824434200, 824435100, 824436000, 824436900, 824437800, 824438700,
    824439600, 824440500, 824441400, 824442300, 824443200, 824444100,
    824445000, 824445900, 824446800, 824447700, 824448600, 824449500,
    824450400, 824451300, 824452200, 824453100, 824454000, 824454900,
    824455800, 824456700, 824457600, 824458500, 824459400, 824460300,
    824461200, 824462100, 824463000, 824463900, 824464800, 824465700,
    824466600, 824467500, 824468400, 824469300, 824470200, 824471100,
    824472000, 824472900, 824473800, 824474700, 824475600, 824476500,
    824477400, 824478300, 824479200, 824480100, 824481000, 824481900,
    824482800, 824483700, 824484600, 824485500, 824486400, 824487300,
    824488200, 824489100, 824490000, 824490900, 824491800, 824492700,
    824493600, 824494500, 824495400, 824496300, 824497200, 824498100,
    824499000, 824499900, 824500800, 824501700, 824502600, 824503500,
    824504400, 824505300, 824506200, 824507100, 824508000, 824508900,
    824509800, 824510700, 824511600, 824512500, 824513400, 824514300,
    824515200, 824516100, 824517000, 824517900, 824518800, 824519700,
    824520600, 824521500, 824522400, 824523300, 824524200, 824525100,
    824526000, 824526900, 824527800, 824528700, 824529600, 824530500,
    824531400, 824532300, 824533200, 824534100, 824535000, 824535900,
    824536800, 824537700, 824538600, 824539500, 824540400, 824541300,
    824542200, 824543100, 824544000, 824544900, 824545800, 824546700,
    824547600, 824548500, 824549400, 824550300, 824551200, 824552100,
    824553000, 824553900, 824554800, 824555700, 824556600, 824557500,
    824558400, 824559300, 824560200, 824561100, 824562000, 824562900,
    824563800, 824564700, 824565600, 824566500, 824567400, 824568300,
    824569200, 824570100, 824571000, 824571900, 824572800, 824573700,
    824574600, 824575500, 824576400, 824577300, 824578200, 824579100,
    824580000, 824580900, 824581800, 824582700, 824583600, 824584500,
    824585400, 824586300, 824587200, 824588100, 824589000, 824589900,
    824590800, 824591700, 824592600, 824593500, 824594400, 824595300,
    824596200, 824597100, 824598000, 824598900, 824599800, 824600700,
    824601600, 824602500, 824603400, 824604300, 824605200, 824606100,
    824607000, 824607900, 824608800, 824609700, 824610600, 824611500,
    824612400, 824613300, 824614200, 824615100, 824616000, 824616900,
    824617800, 824618700, 824619600, 824620500, 824621400, 824622300,
    824623200, 824624100, 824625000, 824625900, 824626800, 824627700,
    824628600, 824629500, 824630400, 824631300, 824632200, 824633100,
    824634000, 824634900, 824635800, 824636700, 824637600, 824638500,
    824639400, 824640300, 824641200, 824642100, 824643000, 824643900,
    824644800, 824645700, 824646600, 824647500, 824648400, 824649300,
    824650200, 824651100, 824652000, 824652900, 824653800, 824654700,
    824655600, 824656500, 824657400, 824658300, 824659200, 824660100,
    824661000, 824661900, 824662800, 824663700, 824664600, 824665500,
    824666400, 824667300, 824668200, 824669100, 824670000, 824670900,
    824671800, 824672700, 824673600, 824674500, 824675400, 824676300,
    824677200, 824678100, 824679000, 824679900, 824680800, 824681700,
    824682600, 824683500, 824684400, 824685300, 824686200, 824687100,
    824688000, 824688900, 824689800, 824690700, 824691600, 824692500,
    824693400, 824694300, 824695200, 824696100, 824697000, 824697900,
    824698800, 824699700, 824700600, 824701500, 824702400, 824703300,
    824704200, 824705100, 824706000, 824706900, 824707800, 824708700,
    824709600, 824710500, 824711400, 824712300, 824713200, 824714100,
    824715000, 824715900, 824716800, 824717700, 824718600, 824719500,
    824720400, 824721300, 824722200, 824723100, 824724000, 824724900,
    824725800, 824726700, 824727600, 824728500, 824729400, 824730300,
    824731200, 824732100, 824733000, 824733900, 824734800, 824735700,
    824736600, 824737500, 824738400, 824739300, 824740200, 824741100,
    824742000, 824742900, 824743800, 824744700, 824745600, 824746500,
    824747400, 824748300, 824749200, 824750100, 824751000, 824751900,
    824752800, 824753700, 824754600, 824755500, 824756400, 824757300,
    824758200, 824759100, 824760000, 824760900, 824761800, 824762700,
    824763600, 824764500, 824765400, 824766300, 824767200, 824768100,
    824769000, 824769900, 824770800, 824771700, 824772600, 824773500,
    824774400, 824775300, 824776200, 824777100, 824778000, 824778900,
    824779800, 824780700, 824781600, 824782500, 824783400, 824784300,
    824785200, 824786100, 824787000, 824787900, 824788800, 824789700,
    824790600, 824791500, 824792400, 824793300, 824794200, 824795100,
    824796000, 824796900, 824797800, 824798700, 824799600, 824800500,
    824801400, 824802300, 824803200, 824804100, 824805000, 824805900,
    824806800, 824807700, 824808600, 824809500, 824810400, 824811300,
    824812200, 824813100, 824814000, 824814900, 824815800, 824816700,
    824817600, 824818500, 824819400, 824820300, 824821200, 824822100,
    824823000, 824823900, 824824800, 824825700, 824826600, 824827500,
    824828400, 824829300, 824830200, 824831100, 824832000, 824832900,
    824833800, 824834700, 824835600, 824836500, 824837400, 824838300,
    824839200, 824840100, 824841000, 824841900, 824842800, 824843700,
    824844600, 824845500, 824846400, 824847300, 824848200, 824849100,
    824850000, 824850900, 824851800, 824852700, 824853600, 824854500,
    824855400, 824856300, 824857200, 824858100, 824859000, 824859900,
    824860800, 824861700, 824862600, 824863500, 824864400, 824865300,
    824866200, 824867100, 824868000, 824868900, 824869800, 824870700,
    824871600, 824872500, 824873400, 824874300, 824875200, 824876100,
    824877000, 824877900, 824878800, 824879700, 824880600, 824881500,
    824882400, 824883300, 824884200, 824885100, 824886000, 824886900,
    824887800, 824888700, 824889600, 824890500, 824891400, 824892300,
    824893200, 824894100, 824895000, 824895900, 824896800, 824897700,
    824898600, 824899500, 824900400, 824901300, 824902200, 824903100,
    824904000, 824904900, 824905800, 824906700, 824907600, 824908500,
    824909400, 824910300, 824911200, 824912100, 824913000, 824913900,
    824914800, 824915700, 824916600, 824917500, 824918400, 824919300,
    824920200, 824921100, 824922000, 824922900, 824923800, 824924700,
    824925600, 824926500, 824927400, 824928300, 824929200, 824930100,
    824931000, 824931900, 824932800, 824933700, 824934600, 824935500,
    824936400, 824937300, 824938200, 824939100, 824940000, 824940900,
    824941800, 824942700, 824943600, 824944500, 824945400, 824946300,
    824947200, 824948100, 824949000, 824949900, 824950800, 824951700,
    824952600, 824953500, 824954400, 824955300, 824956200, 824957100,
    824958000, 824958900, 824959800, 824960700, 824961600, 824962500,
    824963400, 824964300, 824965200, 824966100, 824967000, 824967900,
    824968800, 824969700, 824970600, 824971500, 824972400, 824973300,
    824974200, 824975100, 824976000, 824976900, 824977800, 824978700,
    824979600, 824980500, 824981400, 824982300, 824983200, 824984100,
    824985000, 824985900, 824986800, 824987700, 824988600, 824989500,
    824990400, 824991300, 824992200, 824993100, 824994000, 824994900,
    824995800, 824996700, 824997600, 824998500, 824999400, 825000300,
    825001200, 825002100, 825003000, 825003900, 825004800, 825005700,
    825006600, 825007500, 825008400, 825009300, 825010200, 825011100,
    825012000, 825012900, 825013800, 825014700, 825015600, 825016500,
    825017400, 825018300, 825019200, 825020100, 825021000, 825021900,
    825022800, 825023700, 825024600, 825025500, 825026400, 825027300,
    825028200, 825029100, 825030000, 825030900, 825031800, 825032700,
    825033600, 825034500, 825035400, 825036300, 825037200, 825038100,
    825039000, 825039900, 825040800, 825041700, 825042600, 825043500,
    825044400, 825045300, 825046200, 825047100, 825048000, 825048900,
    825049800, 825050700, 825051600, 825052500, 825053400, 825054300,
    825055200, 825056100, 825057000, 825057900, 825058800, 825059700,
    825060600, 825061500, 825062400, 825063300, 825064200, 825065100,
    825066000, 825066900, 825067800, 825068700, 825069600, 825070500,
    825071400, 825072300, 825073200, 825074100, 825075000, 825075900,
    825076800, 825077700, 825078600, 825079500, 825080400, 825081300,
    825082200, 825083100, 825084000, 825084900, 825085800, 825086700,
    825087600, 825088500, 825089400, 825090300, 825091200, 825092100,
    825093000, 825093900, 825094800, 825095700, 825096600, 825097500,
    825098400, 825099300, 825100200, 825101100, 825102000, 825102900,
    825103800, 825104700, 825105600, 825106500, 825107400, 825108300,
    825109200, 825110100, 825111000, 825111900, 825112800, 825113700,
    825114600, 825115500, 825116400, 825117300, 825118200, 825119100,
    825120000, 825120900, 825121800, 825122700, 825123600, 825124500,
    825125400, 825126300, 825127200, 825128100, 825129000, 825129900,
    825130800, 825131700, 825132600, 825133500, 825134400, 825135300,
    825136200, 825137100, 825138000, 825138900, 825139800, 825140700,
    825141600, 825142500, 825143400, 825144300, 825145200, 825146100,
    825147000, 825147900, 825148800, 825149700, 825150600, 825151500,
    825152400, 825153300, 825154200, 825155100, 825156000, 825156900,
    825157800, 825158700, 825159600, 825160500, 825161400, 825162300,
    825163200, 825164100, 825165000, 825165900, 825166800, 825167700,
    825168600, 825169500, 825170400, 825171300, 825172200, 825173100,
    825174000, 825174900, 825175800, 825176700, 825177600, 825178500,
    825179400, 825180300, 825181200, 825182100, 825183000, 825183900,
    825184800, 825185700, 825186600, 825187500, 825188400, 825189300,
    825190200, 825191100, 825192000, 825192900, 825193800, 825194700,
    825195600, 825196500, 825197400, 825198300, 825199200, 825200100,
    825201000, 825201900, 825202800, 825203700, 825204600, 825205500,
    825206400, 825207300, 825208200, 825209100, 825210000, 825210900,
    825211800, 825212700, 825213600, 825214500, 825215400, 825216300,
    825217200, 825218100, 825219000, 825219900, 825220800, 825221700,
    825222600, 825223500, 825224400, 825225300, 825226200, 825227100,
    825228000, 825228900, 825229800, 825230700, 825231600, 825232500,
    825233400, 825234300, 825235200, 825236100, 825237000, 825237900,
    825238800, 825239700, 825240600, 825241500, 825242400, 825243300,
    825244200, 825245100, 825246000, 825246900, 825247800, 825248700,
    825249600, 825250500, 825251400, 825252300, 825253200, 825254100,
    825255000, 825255900, 825256800, 825257700, 825258600, 825259500,
    825260400, 825261300, 825262200, 825263100, 825264000, 825264900,
    825265800, 825266700, 825267600, 825268500, 825269400, 825270300,
    825271200, 825272100, 825273000, 825273900, 825274800, 825275700,
    825276600, 825277500, 825278400, 825279300, 825280200, 825281100,
    825282000, 825282900, 825283800, 825287400, 825288300, 825289200,
    825290100, 825291000, 825291900, 825292800, 825293700, 825294600,
    825295500, 825296400, 825297300, 825298200, 825299100, 825300000,
    825300900, 825301800, 825302700, 825303600, 825304500, 825305400,
    825306300, 825307200, 825308100, 825309000, 825309900, 825310800,
    825311700, 825312600, 825313500, 825314400, 825315300, 825316200,
    825317100, 825318000, 825318900, 825319800, 825320700, 825321600,
    825322500, 825323400, 825324300, 825325200, 825326100, 825327000,
    825327900, 825328800, 825329700, 825330600, 825331500, 825332400,
    825333300, 825334200, 825335100, 825336000, 825336900, 825337800,
    825338700, 825339600, 825340500, 825341400, 825342300, 825343200,
    825344100, 825345000, 825345900, 825346800, 825347700, 825348600,
    825349500, 825350400, 825351300, 825352200, 825353100, 825354000,
    825354900, 825355800, 825356700, 825357600, 825358500, 825359400,
    825360300, 825361200, 825362100, 825363000, 825363900, 825364800,
    825365700, 825366600, 825367500, 825368400, 825369300, 825370200,
    825371100, 825372000, 825372900, 825373800, 825374700, 825375600,
    825376500, 825377400, 825378300, 825379200, 825380100, 825381000,
    825381900, 825382800, 825383700, 825384600, 825385500, 825386400,
    825387300, 825388200, 825389100, 825390000, 825390900, 825391800,
    825392700, 825393600, 825394500, 825395400, 825396300, 825397200,
    825398100, 825399000, 825399900, 825400800, 825401700, 825402600,
    825403500, 825404400, 825405300, 825406200, 825407100, 825408000,
    825408900, 825409800, 825410700, 825411600, 825412500, 825413400,
    825414300, 825415200, 825416100, 825417000, 825417900, 825418800,
    825419700, 825420600, 825421500, 825422400, 825423300, 825424200,
    825425100, 825426000, 825426900, 825427800, 825428700, 825429600,
    825430500, 825431400, 825432300, 825433200, 825434100, 825435000,
    825435900, 825436800, 825437700, 825438600, 825439500, 825440400,
    825441300, 825442200, 825443100, 825444000, 825444900, 825445800,
    825446700, 825447600, 825448500, 825449400, 825450300, 825451200,
    825452100, 825453000, 825453900, 825454800, 825455700, 825456600,
    825457500, 825458400, 825459300, 825460200, 825461100, 825462000,
    825462900, 825463800, 825464700, 825465600, 825466500, 825467400,
    825468300, 825469200, 825470100, 825471000, 825471900, 825472800,
    825473700, 825474600, 825475500, 825476400, 825477300, 825478200,
    825479100, 825480000, 825480900, 825481800, 825482700, 825483600,
    825484500, 825485400, 825486300, 825487200, 825488100, 825489000,
    825489900, 825490800, 825491700, 825492600, 825493500, 825494400,
    825495300, 825496200, 825497100, 825498000, 825498900, 825499800,
    825500700, 825501600, 825502500, 825503400, 825504300, 825505200,
    825506100, 825507000, 825507900, 825508800, 825509700, 825510600,
    825511500, 825512400, 825513300, 825514200, 825515100, 825516000,
    825516900, 825517800, 825518700, 825519600, 825520500, 825521400,
    825522300, 825523200, 825524100, 825525000, 825525900, 825526800,
    825527700, 825528600, 825529500, 825530400, 825531300, 825532200,
    825533100, 825534000, 825534900, 825535800, 825536700, 825537600,
    825538500, 825539400, 825540300, 825541200, 825542100, 825543000,
    825543900, 825544800, 825545700, 825546600, 825547500, 825548400,
    825549300, 825550200, 825551100, 825552000, 825552900, 825553800,
    825554700, 825555600, 825556500, 825557400, 825558300, 825559200,
    825560100, 825561000, 825561900, 825562800, 825563700, 825564600,
    825565500, 825566400, 825567300, 825568200, 825569100, 825570000,
    825570900, 825571800, 825572700, 825573600, 825574500, 825575400,
    825576300, 825577200, 825578100, 825579000, 825579900, 825580800,
    825581700, 825582600, 825583500, 825584400, 825585300, 825586200,
    825587100, 825588000, 825588900, 825589800, 825590700, 825591600,
    825592500, 825593400, 825594300, 825595200, 825596100, 825597000,
    825597900, 825598800, 825599700, 825600600, 825601500, 825602400,
    825603300, 825604200, 825605100, 825606000, 825606900, 825607800,
    825608700, 825609600, 825610500, 825611400, 825612300, 825613200,
    825614100, 825615000, 825615900, 825616800, 825617700, 825618600,
    825619500, 825620400, 825621300, 825622200, 825623100, 825624000,
    825624900, 825625800, 825626700, 825627600, 825628500, 825629400,
    825630300, 825631200, 825632100, 825633000, 825633900, 825634800,
    825635700, 825636600, 825637500, 825638400, 825639300, 825640200,
    825641100, 825642000, 825642900, 825643800, 825644700, 825645600,
    825646500, 825647400, 825648300, 825649200, 825650100, 825651000,
    825651900, 825652800, 825653700, 825654600, 825655500, 825656400,
    825657300, 825658200, 825659100, 825660000, 825660900, 825661800,
    825662700, 825663600, 825664500, 825665400, 825666300, 825667200,
    825668100, 825669000, 825669900, 825670800, 825671700, 825672600,
    825673500, 825674400, 825675300, 825676200, 825677100, 825678000,
    825678900, 825679800, 825680700, 825681600, 825682500, 825683400,
    825684300, 825685200, 825686100, 825687000, 825687900, 825688800,
    825689700, 825690600, 825691500, 825692400, 825693300, 825694200,
    825695100, 825696000, 825696900, 825697800, 825698700, 825699600,
    825700500, 825701400, 825702300, 825703200, 825704100, 825705000,
    825705900, 825706800, 825707700, 825708600, 825709500, 825710400,
    825711300, 825712200, 825713100, 825714000, 825714900, 825715800,
    825716700, 825717600, 825718500, 825719400, 825720300, 825721200,
    825722100, 825723000, 825723900, 825724800, 825725700, 825726600,
    825727500, 825728400, 825729300, 825730200, 825731100, 825732000,
    825732900, 825733800, 825734700, 825735600, 825736500, 825737400,
    825738300, 825739200, 825740100, 825741000, 825741900, 825742800,
    825743700, 825744600, 825745500, 825746400, 825747300, 825748200,
    825749100, 825750000, 825750900, 825751800, 825752700, 825753600,
    825754500, 825755400, 825756300, 825757200, 825758100, 825759000,
    825759900, 825760800, 825761700, 825762600, 825763500, 825764400,
    825765300, 825766200, 825767100, 825768000, 825768900, 825769800,
    825770700, 825771600, 825772500, 825773400, 825774300, 825775200,
    825776100, 825777000, 825777900, 825778800, 825779700, 825780600,
    825781500, 825782400, 825783300, 825784200, 825785100, 825786000,
    825786900, 825787800, 825788700, 825789600, 825790500, 825791400,
    825792300, 825793200, 825794100, 825795000, 825795900, 825796800,
    825797700, 825798600, 825799500, 825800400, 825801300, 825802200,
    825803100, 825804000, 825804900, 825805800, 825806700, 825807600,
    825808500, 825809400, 825810300, 825811200, 825812100, 825813000,
    825813900, 825814800, 825815700, 825816600, 825817500, 825818400,
    825819300, 825820200, 825821100, 825822000, 825822900, 825823800,
    825824700, 825825600, 825826500, 825827400, 825828300, 825829200,
    825830100, 825831000, 825831900, 825832800, 825833700, 825834600,
    825835500, 825836400, 825837300, 825838200, 825839100, 825840000,
    825840900, 825841800, 825842700, 825843600, 825844500, 825845400,
    825846300, 825847200, 825848100, 825849000, 825849900, 825850800,
    825851700, 825852600, 825853500, 825854400, 825855300, 825856200,
    825857100, 825858000, 825858900, 825859800, 825860700, 825861600,
    825862500, 825863400, 825864300, 825865200, 825866100, 825867000,
    825867900, 825868800, 825869700, 825870600, 825871500, 825872400,
    825873300, 825874200, 825875100, 825876000, 825876900, 825877800,
    825878700, 825879600, 825880500, 825881400, 825882300, 825883200,
    825884100, 825885000, 825885900, 825886800, 825887700, 825888600,
    825889500, 825890400, 825891300, 825892200, 825893100, 825894000,
    825894900, 825895800, 825896700, 825897600, 825898500, 825899400,
    825900300, 825901200, 825902100, 825903000, 825903900, 825904800,
    825905700, 825906600, 825907500, 825908400, 825909300, 825910200,
    825911100, 825912000, 825912900, 825913800, 825914700, 825915600,
    825916500, 825917400, 825918300, 825919200, 825920100, 825921000,
    825921900, 825922800, 825923700, 825924600, 825925500, 825926400,
    825927300, 825928200, 825929100, 825930000, 825930900, 825931800,
    825932700, 825933600, 825934500, 825935400, 825936300, 825937200,
    825938100, 825939000, 825939900, 825940800, 825941700, 825942600,
    825943500, 825944400, 825945300, 825946200, 825947100, 825948000,
    825948900, 825949800, 825950700, 825951600, 825952500, 825953400,
    825954300, 825955200, 825956100, 825957000, 825957900, 825958800,
    825959700, 825960600, 825961500, 825962400, 825963300, 825964200,
    825965100, 825966000, 825966900, 825967800, 825968700, 825969600,
    825970500, 825971400, 825972300, 825973200, 825974100, 825975000,
    825975900, 825976800, 825977700, 825978600, 825979500, 825980400,
    825981300, 825982200, 825983100, 825984000, 825984900, 825985800,
    825986700, 825987600, 825988500, 825989400, 825990300, 825991200,
    825992100, 825993000, 825993900, 825994800, 825995700, 825996600,
    825997500, 825998400, 825999300, 826000200, 826001100, 826002000,
    826002900, 826003800, 826004700, 826005600, 826006500, 826007400,
    826008300, 826009200, 826010100, 826011000, 826011900, 826012800,
    826013700, 826014600, 826015500, 826016400, 826017300, 826018200,
    826019100, 826020000, 826020900, 826021800, 826022700, 826023600,
    826024500, 826025400, 826026300, 826027200, 826028100, 826029000,
    826029900, 826030800, 826031700, 826032600, 826033500, 826034400,
    826035300, 826036200, 826037100, 826038000, 826038900, 826039800,
    826040700, 826041600, 826042500, 826043400, 826044300, 826045200,
    826046100, 826047000, 826047900, 826048800, 826049700, 826050600,
    826051500, 826052400, 826053300, 826054200, 826055100, 826056000,
    826056900, 826057800, 826058700, 826059600, 826060500, 826061400,
    826062300, 826063200, 826064100, 826065000, 826065900, 826066800,
    826067700, 826068600, 826069500, 826070400, 826071300, 826072200,
    826073100, 826074000, 826074900, 826075800, 826076700, 826077600,
    826078500, 826079400, 826080300, 826081200, 826082100, 826083000,
    826083900, 826084800, 826085700, 826086600, 826087500, 826088400,
    826089300, 826090200, 826091100, 826092000, 826092900, 826093800,
    826094700, 826095600, 826096500, 826097400, 826098300, 826099200,
    826100100, 826101000, 826101900, 826102800, 826103700, 826104600,
    826105500, 826106400, 826107300, 826108200, 826109100, 826110000,
    826110900, 826111800, 826112700, 826113600, 826114500, 826115400,
    826116300, 826117200, 826118100, 826119000, 826119900, 826120800,
    826121700, 826122600, 826123500, 826124400, 826125300, 826126200,
    826127100, 826128000, 826128900, 826129800, 826130700, 826131600,
    826132500, 826133400, 826134300, 826135200, 826136100, 826137000,
    826137900, 826138800, 826139700, 826140600, 826141500, 826142400,
    826143300, 826144200, 826145100, 826146000, 826146900, 826147800,
    826148700, 826149600, 826150500, 826151400, 826152300, 826153200,
    826154100, 826155000, 826155900, 826156800, 826157700, 826158600,
    826159500, 826160400, 826161300, 826162200, 826163100, 826164000,
    826164900, 826165800, 826166700, 826167600, 826168500, 826169400,
    826170300, 826171200, 826172100, 826173000, 826173900, 826174800,
    826175700, 826176600, 826177500, 826178400, 826179300, 826180200,
    826181100, 826182000, 826182900, 826183800, 826184700, 826185600,
    826186500, 826187400, 826188300, 826189200, 826190100, 826191000,
    826191900, 826192800, 826193700, 826194600, 826195500, 826196400,
    826197300, 826198200, 826199100, 826200000, 826200900, 826201800,
    826202700, 826203600, 826204500, 826205400, 826206300, 826207200,
    826208100, 826209000, 826209900, 826210800, 826211700, 826212600,
    826213500, 826214400, 826215300, 826216200, 826217100, 826218000,
    826218900, 826219800, 826220700, 826221600, 826222500, 826223400,
    826224300, 826225200, 826226100, 826227000, 826227900, 826228800,
    826229700, 826230600, 826231500, 826232400, 826233300, 826234200,
    826235100, 826236000, 826236900, 826237800, 826238700, 826239600,
    826240500, 826241400, 826242300, 826243200, 826244100, 826245000,
    826245900, 826246800, 826247700, 826248600, 826249500, 826250400,
    826251300, 826252200, 826253100, 826254000, 826254900, 826255800,
    826256700, 826257600, 826258500, 826259400, 826260300, 826261200,
    826262100, 826263000, 826263900, 826264800, 826265700, 826266600,
    826267500, 826268400, 826269300, 826270200, 826271100, 826272000,
    826272900, 826273800, 826274700, 826275600, 826276500, 826277400,
    826278300, 826279200, 826280100, 826281000, 826281900, 826282800,
    826283700, 826284600, 826285500, 826286400, 826287300, 826288200,
    826289100, 826290000, 826290900, 826291800, 826292700, 826293600,
    826294500, 826295400, 826296300, 826297200, 826298100, 826299000,
    826299900, 826300800, 826301700, 826302600, 826303500, 826304400,
    826305300, 826306200, 826307100, 826308000, 826308900, 826309800,
    826310700, 826311600, 826312500, 826313400, 826314300, 826315200,
    826316100, 826317000, 826317900, 826318800, 826319700, 826320600,
    826321500, 826322400, 826323300, 826324200, 826325100, 826326000,
    826326900, 826327800, 826328700, 826329600, 826330500, 826331400,
    826332300, 826333200, 826334100, 826335000, 826335900, 826336800,
    826337700, 826338600, 826339500, 826340400, 826341300, 826342200,
    826343100, 826344000, 826344900, 826345800, 826346700, 826347600,
    826348500, 826349400, 826350300, 826351200, 826352100, 826353000,
    826353900, 826354800, 826355700, 826356600, 826357500, 826358400,
    826359300, 826360200, 826361100, 826362000, 826362900, 826363800,
    826364700, 826365600, 826366500, 826367400, 826368300, 826369200,
    826370100, 826371000, 826371900, 826372800, 826373700, 826374600,
    826375500, 826376400, 826377300, 826378200, 826379100, 826380000,
    826380900, 826381800, 826382700, 826383600, 826384500, 826385400,
    826386300, 826387200, 826388100, 826389000, 826389900, 826390800,
    826391700, 826392600, 826393500, 826394400, 826395300, 826396200,
    826397100, 826398000, 826398900, 826399800, 826400700, 826401600,
    826402500, 826403400, 826404300, 826405200, 826406100, 826407000,
    826407900, 826408800, 826409700, 826410600, 826411500, 826412400,
    826413300, 826414200, 826415100, 826416000, 826416900, 826417800,
    826418700, 826419600, 826420500, 826421400, 826422300, 826423200,
    826424100, 826425000, 826425900, 826426800, 826427700, 826428600,
    826429500, 826430400, 826431300, 826432200, 826433100, 826434000,
    826434900, 826435800, 826436700, 826437600, 826438500, 826439400,
    826440300, 826441200, 826442100, 826443000, 826443900, 826444800,
    826445700, 826446600, 826447500, 826448400, 826449300, 826450200,
    826451100, 826452000, 826452900, 826453800, 826454700, 826455600,
    826456500, 826457400, 826458300, 826459200, 826460100, 826461000,
    826461900, 826462800, 826463700, 826464600, 826465500, 826466400,
    826467300, 826468200, 826469100, 826470000, 826470900, 826471800,
    826472700, 826473600, 826474500, 826475400, 826476300, 826477200,
    826478100, 826479000, 826479900, 826480800, 826481700, 826482600,
    826483500, 826484400, 826485300, 826486200, 826487100, 826488000,
    826488900, 826489800, 826490700, 826491600, 826492500, 826493400,
    826494300, 826495200, 826496100, 826497000, 826497900, 826498800,
    826499700, 826500600, 826501500, 826502400, 826503300, 826504200,
    826505100, 826506000, 826506900, 826507800, 826508700, 826509600,
    826510500, 826511400, 826512300, 826513200, 826514100, 826515000,
    826515900, 826516800, 826517700, 826518600, 826519500, 826520400,
    826521300, 826522200, 826523100, 826524000, 826524900, 826525800,
    826526700, 826527600, 826528500, 826529400, 826530300, 826531200,
    826532100, 826533000, 826533900, 826534800, 826535700, 826536600,
    826537500, 826538400, 826539300, 826540200, 826541100, 826542000,
    826542900, 826543800, 826544700, 826545600, 826546500, 826547400,
    826548300, 826549200, 826550100, 826551000, 826551900, 826552800,
    826553700, 826554600, 826555500, 826556400, 826557300, 826558200,
    826559100, 826560000, 826560900, 826561800, 826562700, 826563600,
    826564500, 826565400, 826566300, 826567200, 826568100, 826569000,
    826569900, 826570800, 826571700, 826572600, 826573500, 826574400,
    826575300, 826576200, 826577100, 826578000, 826578900, 826579800,
    826580700, 826581600, 826582500, 826583400, 826584300, 826585200,
    826586100, 826587000, 826587900, 826588800, 826589700, 826590600,
    826591500, 826592400, 826593300, 826594200, 826595100, 826596000,
    826596900, 826597800, 826598700, 826599600, 826600500, 826601400,
    826602300, 826603200, 826604100, 826605000, 826605900, 826606800,
    826607700, 826608600, 826609500, 826610400, 826611300, 826612200,
    826613100, 826614000, 826614900, 826615800, 826616700, 826617600,
    826618500, 826619400, 826620300, 826621200, 826622100, 826623000,
    826623900, 826624800, 826625700, 826626600, 826627500, 826628400,
    826629300, 826630200, 826631100, 826632000, 826632900, 826633800,
    826634700, 826635600, 826636500, 826637400, 826638300, 826639200,
    826640100, 826641000, 826641900, 826642800, 826643700, 826644600,
    826645500, 826646400, 826647300, 826648200, 826649100, 826650000,
    826650900, 826651800, 826652700, 826653600, 826654500, 826655400,
    826656300, 826657200, 826658100, 826659000, 826659900, 826660800,
    826661700, 826662600, 826663500, 826664400, 826665300, 826666200,
    826667100, 826668000, 826668900, 826669800, 826670700, 826671600,
    826672500, 826673400, 826674300, 826675200, 826676100, 826677000,
    826677900, 826678800, 826679700, 826680600, 826681500, 826682400,
    826683300, 826684200, 826685100, 826686000, 826686900, 826687800,
    826688700, 826689600, 826690500, 826691400, 826692300, 826693200,
    826694100, 826695000, 826695900, 826696800, 826697700, 826698600,
    826699500, 826700400, 826701300, 826702200, 826703100, 826704000,
    826704900, 826705800, 826706700, 826707600, 826708500, 826709400,
    826710300, 826711200, 826712100, 826713000, 826713900, 826714800,
    826715700, 826716600, 826717500, 826718400, 826719300, 826720200,
    826721100, 826722000, 826722900, 826723800, 826724700, 826725600,
    826726500, 826727400, 826728300, 826729200, 826730100, 826731000,
    826731900, 826732800, 826733700, 826734600, 826735500, 826736400,
    826737300, 826738200, 826739100, 826740000, 826740900, 826741800,
    826742700, 826743600, 826744500, 826745400, 826746300, 826747200,
    826748100, 826749000, 826749900, 826750800, 826751700, 826752600,
    826753500, 826754400, 826755300, 826756200, 826757100, 826758000,
    826758900, 826759800, 826760700, 826761600, 826762500, 826763400,
    826764300, 826765200, 826766100, 826767000, 826767900, 826768800,
    826769700, 826770600, 826771500, 826772400, 826773300, 826774200,
    826775100, 826776000, 826776900, 826777800, 826778700, 826779600,
    826780500, 826781400, 826782300, 826783200, 826784100, 826785000,
    826785900, 826786800, 826787700, 826788600, 826789500, 826790400,
    826791300, 826792200, 826793100, 826794000, 826794900, 826795800,
    826796700, 826797600, 826798500, 826799400, 826800300, 826801200,
    826802100, 826803000, 826803900, 826804800, 826805700, 826806600,
    826807500, 826808400, 826809300, 826810200, 826811100, 826812000,
    826812900, 826813800, 826814700, 826815600, 826816500, 826817400,
    826818300, 826819200, 826820100, 826821000, 826821900, 826822800,
    826823700, 826824600, 826825500, 826826400, 826827300, 826828200,
    826829100, 826830000, 826830900, 826831800, 826832700, 826833600,
    826834500, 826835400, 826836300, 826837200, 826838100, 826839000,
    826839900, 826840800, 826841700, 826842600, 826843500, 826844400,
    826845300, 826846200, 826847100, 826848000, 826848900, 826849800,
    826850700, 826851600, 826852500, 826853400, 826854300, 826855200,
    826856100, 826857000, 826857900, 826858800, 826859700, 826860600,
    826861500, 826862400, 826863300, 826864200, 826865100, 826866000,
    826866900, 826867800, 826868700, 826869600, 826870500, 826871400,
    826872300, 826873200, 826874100, 826875000, 826875900, 826876800,
    826877700, 826878600, 826879500, 826880400, 826881300, 826882200,
    826883100, 826884000, 826884900, 826885800, 826886700, 826887600,
    826888500, 826889400, 826890300, 826891200, 826892100, 826893000,
    826893900, 826894800, 826895700, 826896600, 826897500, 826898400,
    826899300, 826900200, 826901100, 826902000, 826902900, 826903800,
    826904700, 826905600, 826906500, 826907400, 826908300, 826909200,
    826910100, 826911000, 826911900, 826912800, 826913700, 826914600,
    826915500, 826916400, 826917300, 826918200, 826919100, 826920000,
    826920900, 826921800, 826922700, 826923600, 826924500, 826925400,
    826926300, 826927200, 826928100, 826929000, 826929900, 826930800,
    826931700, 826932600, 826933500, 826934400, 826935300, 826936200,
    826937100, 826938000, 826938900, 826939800, 826940700, 826941600,
    826942500, 826943400, 826944300, 826945200, 826946100, 826947000,
    826947900, 826948800, 826949700, 826950600, 826951500, 826952400,
    826953300, 826954200, 826955100, 826956000, 826956900, 826957800,
    826958700, 826959600, 826960500, 826961400, 826962300, 826963200,
    826964100, 826965000, 826965900, 826966800, 826967700, 826968600,
    826969500, 826970400, 826971300, 826972200, 826973100, 826974000,
    826974900, 826975800, 826976700, 826977600, 826978500, 826979400,
    826980300, 826981200, 826982100, 826983000, 826983900, 826984800,
    826985700, 826986600, 826987500, 826988400, 826989300, 826990200,
    826991100, 826992000, 826992900, 826993800, 826994700, 826995600,
    826996500, 826997400, 826998300, 826999200, 827000100, 827001000,
    827001900, 827002800, 827003700, 827004600, 827005500, 827006400,
    827007300, 827008200, 827009100, 827010000, 827010900, 827011800,
    827012700, 827013600, 827014500, 827015400, 827016300, 827017200,
    827018100, 827019000, 827019900, 827020800, 827021700, 827022600,
    827023500, 827024400, 827025300, 827026200, 827027100, 827028000,
    827028900, 827029800, 827030700, 827031600, 827032500, 827033400,
    827034300, 827035200, 827036100, 827037000, 827037900, 827038800,
    827039700, 827040600, 827041500, 827042400, 827043300, 827044200,
    827045100, 827046000, 827046900, 827047800, 827048700, 827049600,
    827050500, 827051400, 827052300, 827053200, 827054100, 827055000,
    827055900, 827056800, 827057700, 827058600, 827059500, 827060400,
    827061300, 827062200, 827063100, 827064000, 827064900, 827065800,
    827066700, 827067600, 827068500, 827069400, 827070300, 827071200,
    827072100, 827073000, 827073900, 827074800, 827075700, 827076600,
    827077500, 827078400, 827079300, 827080200, 827081100, 827082000,
    827082900, 827083800, 827084700, 827085600, 827086500, 827087400,
    827088300, 827089200, 827090100, 827091000, 827091900, 827092800,
    827093700, 827094600, 827095500, 827096400, 827097300, 827098200,
    827099100, 827100000, 827100900, 827101800, 827102700, 827103600,
    827104500, 827105400, 827106300, 827107200, 827108100, 827109000,
    827109900, 827110800, 827111700, 827112600, 827113500, 827114400,
    827115300, 827116200, 827117100, 827118000, 827118900, 827119800,
    827120700, 827121600, 827122500, 827123400, 827124300, 827125200,
    827126100, 827127000, 827127900, 827128800, 827129700, 827130600,
    827131500, 827132400, 827133300, 827134200, 827135100, 827136000,
    827136900, 827137800, 827138700, 827139600, 827140500, 827141400,
    827142300, 827143200, 827144100, 827145000, 827145900, 827146800,
    827147700, 827148600, 827149500, 827150400, 827151300, 827152200,
    827153100, 827154000, 827154900, 827155800, 827156700, 827157600,
    827158500, 827159400, 827160300, 827161200, 827162100, 827163000,
    827163900, 827164800, 827165700, 827166600, 827167500, 827168400,
    827169300, 827170200, 827171100, 827172000, 827172900, 827173800,
    827174700, 827175600, 827176500, 827177400, 827178300, 827179200,
    827180100, 827181000, 827181900, 827182800, 827183700, 827184600,
    827185500, 827186400, 827187300, 827188200, 827189100, 827190000,
    827190900, 827191800, 827192700, 827193600, 827194500, 827195400,
    827196300, 827197200, 827198100, 827199000, 827199900, 827200800,
    827201700, 827202600, 827203500, 827204400, 827205300, 827206200,
    827207100, 827208000, 827208900, 827209800, 827210700, 827211600,
    827212500, 827213400, 827214300, 827215200, 827216100, 827217000,
    827217900, 827218800, 827219700, 827220600, 827221500, 827222400,
    827223300, 827224200, 827225100, 827226000, 827226900, 827227800,
    827228700, 827229600, 827230500, 827231400, 827232300, 827233200,
    827234100, 827235000, 827235900, 827236800, 827237700, 827238600,
    827239500, 827240400, 827241300, 827242200, 827243100, 827244000,
    827244900, 827245800, 827246700, 827247600, 827248500, 827249400,
    827250300, 827251200, 827252100, 827253000, 827253900, 827254800,
    827255700, 827256600, 827257500, 827258400, 827259300, 827260200,
    827261100, 827262000, 827262900, 827263800, 827264700, 827265600,
    827266500, 827267400, 827268300, 827269200, 827270100, 827271000,
    827271900, 827272800, 827273700, 827274600, 827275500, 827276400,
    827277300, 827278200, 827279100, 827280000, 827280900, 827281800,
    827282700, 827283600, 827284500, 827285400, 827286300, 827287200,
    827288100, 827289000, 827289900, 827290800, 827291700, 827292600,
    827293500, 827294400, 827295300, 827296200, 827297100, 827298000,
    827298900, 827299800, 827300700, 827301600, 827302500, 827303400,
    827304300, 827305200, 827306100, 827307000, 827307900, 827308800,
    827309700, 827310600, 827311500, 827312400, 827313300, 827314200,
    827315100, 827316000, 827316900, 827317800, 827318700, 827319600,
    827320500, 827321400, 827322300, 827323200, 827324100, 827325000,
    827325900, 827326800, 827327700, 827328600, 827329500, 827330400,
    827331300, 827332200, 827333100, 827334000, 827334900, 827335800,
    827336700, 827337600, 827338500, 827339400, 827340300, 827341200,
    827342100, 827343000, 827343900, 827344800, 827345700, 827346600,
    827347500, 827348400, 827349300, 827350200, 827351100, 827352000,
    827352900, 827353800, 827354700, 827355600, 827356500, 827357400,
    827358300, 827359200, 827360100, 827361000, 827361900, 827362800,
    827363700, 827364600, 827365500, 827366400, 827367300, 827368200,
    827369100, 827370000, 827370900, 827371800, 827372700, 827373600,
    827374500, 827375400, 827376300, 827377200, 827378100, 827379000,
    827379900, 827380800, 827381700, 827382600, 827383500, 827384400,
    827385300, 827386200, 827387100, 827388000, 827388900, 827389800,
    827390700, 827391600, 827392500, 827393400, 827394300, 827395200,
    827396100, 827397000, 827397900, 827398800, 827399700, 827400600,
    827401500, 827402400, 827403300, 827404200, 827405100, 827406000,
    827406900, 827407800, 827408700, 827409600, 827410500, 827411400,
    827412300, 827413200, 827414100, 827415000, 827415900, 827416800,
    827417700, 827418600, 827419500, 827420400, 827421300, 827422200,
    827423100, 827424000, 827424900, 827425800, 827426700, 827427600,
    827428500, 827429400, 827430300, 827431200, 827432100, 827433000,
    827433900, 827434800, 827435700, 827436600, 827437500, 827438400,
    827439300, 827440200, 827441100, 827442000, 827442900, 827443800,
    827444700, 827445600, 827446500, 827447400, 827448300, 827449200,
    827450100, 827451000, 827451900, 827452800, 827453700, 827454600,
    827455500, 827456400, 827457300, 827458200, 827459100, 827460000,
    827460900, 827461800, 827462700, 827463600, 827464500, 827465400,
    827466300, 827467200, 827468100, 827469000, 827469900, 827470800,
    827471700, 827472600, 827473500, 827474400, 827475300, 827476200,
    827477100, 827478000, 827478900, 827479800, 827480700, 827481600,
    827482500, 827483400, 827484300, 827485200, 827486100, 827487000,
    827487900, 827488800, 827489700, 827490600, 827491500, 827492400,
    827493300, 827494200, 827495100, 827496000, 827496900, 827497800,
    827498700, 827499600, 827500500, 827501400, 827502300, 827503200,
    827504100, 827505000, 827505900, 827506800, 827507700, 827508600,
    827509500, 827510400, 827511300, 827512200, 827513100, 827514000,
    827514900, 827515800, 827516700, 827517600, 827518500, 827519400,
    827520300, 827521200, 827522100, 827523000, 827523900, 827524800,
    827525700, 827526600, 827527500, 827528400, 827529300, 827530200,
    827531100, 827532000, 827532900, 827533800, 827534700, 827535600,
    827536500, 827537400, 827538300, 827539200, 827540100, 827541000,
    827541900, 827542800, 827543700, 827544600, 827545500, 827546400,
    827547300, 827548200, 827549100, 827550000, 827550900, 827551800,
    827552700, 827553600, 827554500, 827555400, 827556300, 827557200,
    827558100, 827559000, 827559900, 827560800, 827561700, 827562600,
    827563500, 827564400, 827565300, 827566200, 827567100, 827568000,
    827568900, 827569800, 827570700, 827571600, 827572500, 827573400,
    827574300, 827575200, 827576100, 827577000, 827577900, 827578800,
    827579700, 827580600, 827581500, 827582400, 827583300, 827584200,
    827585100, 827586000, 827586900, 827587800, 827588700, 827589600,
    827590500, 827591400, 827592300, 827593200, 827594100, 827595000,
    827595900, 827596800, 827597700, 827598600, 827599500, 827600400,
    827601300, 827602200, 827603100, 827604000, 827604900, 827605800,
    827606700, 827607600, 827608500, 827609400, 827610300, 827611200,
    827612100, 827613000, 827613900, 827614800, 827615700, 827616600,
    827617500, 827618400, 827619300, 827620200, 827621100, 827622000,
    827622900, 827623800, 827624700, 827625600, 827626500, 827627400,
    827628300, 827629200, 827630100, 827631000, 827631900, 827632800,
    827633700, 827634600, 827635500, 827636400, 827637300, 827638200,
    827639100, 827640000, 827640900, 827641800, 827642700, 827643600,
    827644500, 827645400, 827646300, 827647200, 827648100, 827649000,
    827649900, 827650800, 827651700, 827652600, 827653500, 827654400,
    827655300, 827656200, 827657100, 827658000, 827658900, 827659800,
    827660700, 827661600, 827662500, 827663400, 827664300, 827665200,
    827666100, 827667000, 827667900, 827668800, 827669700, 827670600,
    827671500, 827672400, 827673300, 827674200, 827675100, 827676000,
    827676900, 827677800, 827678700, 827679600, 827680500, 827681400,
    827682300, 827683200, 827684100, 827685000, 827685900, 827686800,
    827687700, 827688600, 827689500, 827690400, 827691300, 827692200,
    827693100, 827694000, 827694900, 827695800, 827696700, 827697600,
    827698500, 827699400, 827700300, 827701200, 827702100, 827703000,
    827703900, 827704800, 827705700, 827706600, 827707500, 827708400,
    827709300, 827710200, 827711100, 827712000, 827712900, 827713800,
    827714700, 827715600, 827716500, 827717400, 827718300, 827719200,
    827720100, 827721000, 827721900, 827722800, 827723700, 827724600,
    827725500, 827726400, 827727300, 827728200, 827729100, 827730000,
    827730900, 827731800, 827732700, 827733600, 827734500, 827735400,
    827736300, 827737200, 827738100, 827739000, 827739900, 827740800,
    827741700, 827742600, 827743500, 827744400, 827745300, 827746200,
    827747100, 827748000, 827748900, 827749800, 827750700, 827751600,
    827752500, 827753400, 827754300, 827755200, 827756100, 827757000,
    827757900, 827758800, 827759700, 827760600, 827761500, 827762400,
    827763300, 827764200, 827765100, 827766000, 827766900, 827767800,
    827768700, 827769600, 827770500, 827771400, 827772300, 827773200,
    827774100, 827775000, 827775900, 827776800, 827777700, 827778600,
    827783100, 827784000, 827784900, 827785800, 827786700, 827787600,
    827788500, 827789400, 827790300, 827791200, 827792100, 827793000,
    827793900, 827794800, 827795700, 827796600, 827797500, 827798400,
    827799300, 827800200, 827801100, 827802000, 827802900, 827803800,
    827804700, 827805600, 827806500, 827807400, 827808300, 827809200,
    827810100, 827811000, 827811900, 827812800, 827813700, 827814600,
    827815500, 827816400, 827817300, 827818200, 827819100, 827820000,
    827820900, 827821800, 827822700, 827823600, 827824500, 827825400,
    827826300, 827827200, 827828100, 827829000, 827829900, 827830800,
    827831700, 827832600, 827833500, 827834400, 827835300, 827836200,
    827837100, 827838000, 827838900, 827839800, 827840700, 827841600,
    827842500, 827843400, 827844300, 827845200, 827846100, 827847000,
    827847900, 827848800, 827849700, 827850600, 827851500, 827852400,
    827853300, 827854200, 827855100, 827856000, 827856900, 827857800,
    827858700, 827859600, 827860500, 827861400, 827862300, 827863200,
    827864100, 827865000, 827865900, 827866800, 827867700, 827868600,
    827869500, 827870400, 827871300, 827872200, 827873100, 827874000,
    827874900, 827875800, 827876700, 827877600, 827878500, 827879400,
    827880300, 827881200, 827882100, 827883000, 827883900, 827884800,
    827885700, 827886600, 827887500, 827888400, 827889300, 827890200,
    827891100, 827892000, 827892900, 827893800, 827894700, 827895600,
    827896500, 827897400, 827898300, 827899200, 827900100, 827901000,
    827901900, 827902800, 827903700, 827904600, 827905500, 827906400,
    827907300, 827908200, 827909100, 827910000, 827910900, 827911800,
    827912700, 827913600, 827914500, 827915400, 827916300, 827917200,
    827918100, 827919000, 827919900, 827920800, 827921700, 827922600,
    827923500, 827924400, 827925300, 827926200, 827927100, 827928000,
    827928900, 827929800, 827930700, 827931600, 827932500, 827933400,
    827934300, 827935200, 827936100, 827937000, 827937900, 827938800,
    827939700, 827940600, 827941500, 827942400, 827943300, 827944200,
    827945100, 827946000, 827946900, 827947800, 827948700, 827949600,
    827950500, 827951400, 827952300, 827953200, 827954100, 827955000,
    827955900, 827956800, 827957700, 827958600, 827959500, 827960400,
    827961300, 827962200, 827963100, 827964000, 827964900, 827965800,
    827966700, 827967600, 827968500, 827969400, 827970300, 827971200,
    827972100, 827973000, 827973900, 827974800, 827975700, 827976600,
    827977500, 827978400, 827979300, 827980200, 827981100, 827982000,
    827982900, 827983800, 827984700, 827985600, 827986500, 827987400,
    827988300, 827989200, 827990100, 827991000, 827991900, 827992800,
    827993700, 827994600, 827995500, 827996400, 827997300, 827998200,
    827999100, 828000000, 828000900, 828001800, 828002700, 828003600,
    828004500, 828005400, 828006300, 828007200, 828008100, 828009000,
    828009900, 828010800, 828011700, 828012600, 828013500, 828014400,
    828015300, 828016200, 828017100, 828018000, 828018900, 828019800,
    828020700, 828021600, 828022500, 828023400, 828024300, 828025200,
    828026100, 828027000, 828027900, 828028800, 828029700, 828030600,
    828031500, 828032400, 828033300, 828034200, 828035100, 828036000,
    828036900, 828037800, 828038700, 828039600, 828040500, 828041400,
    828042300, 828043200, 828044100, 828045000, 828045900, 828046800,
    828047700, 828048600, 828049500, 828050400, 828051300, 828052200,
    828053100, 828054000, 828054900, 828055800, 828056700, 828057600,
    828058500, 828059400, 828060300, 828061200, 828062100, 828063000,
    828063900, 828064800, 828065700, 828066600, 828067500, 828068400,
    828069300, 828070200, 828071100, 828072000, 828072900, 828073800,
    828074700, 828075600, 828076500, 828077400, 828078300, 828079200,
    828080100, 828081000, 828081900, 828082800, 828083700, 828084600,
    828085500, 828086400, 828087300, 828088200, 828089100, 828090000,
    828090900, 828091800, 828092700, 828093600, 828094500, 828095400,
    828096300, 828097200, 828098100, 828099000, 828099900, 828100800,
    828101700, 828102600, 828103500, 828104400, 828105300, 828106200,
    828107100, 828108000, 828108900, 828109800, 828110700, 828111600,
    828112500, 828113400, 828114300, 828115200, 828116100, 828117000,
    828117900, 828118800, 828119700, 828120600, 828121500, 828122400,
    828123300, 828124200, 828125100, 828126000, 828126900, 828127800,
    828128700, 828129600, 828130500, 828131400, 828132300, 828133200,
    828134100, 828135000, 828135900, 828136800, 828137700, 828138600,
    828139500, 828140400, 828141300, 828142200, 828143100, 828144000,
    828144900, 828145800, 828146700, 828147600, 828148500, 828149400,
    828150300, 828151200, 828152100, 828153000, 828153900, 828154800,
    828155700, 828156600, 828157500, 828158400, 828159300, 828160200,
    828161100, 828162000, 828162900, 828163800, 828164700, 828165600,
    828166500, 828167400, 828168300, 828169200, 828170100, 828171000,
    828171900, 828172800, 828173700, 828174600, 828175500, 828176400,
    828177300, 828178200, 828179100, 828180000, 828180900, 828181800,
    828182700, 828183600, 828184500, 828185400, 828186300, 828187200,
    828188100, 828189000, 828189900, 828190800, 828191700, 828192600,
    828193500, 828194400, 828195300, 828196200, 828197100, 828198000,
    828198900, 828199800, 828200700, 828201600, 828202500, 828203400,
    828204300, 828205200, 828206100, 828207000, 828207900, 828208800,
    828209700, 828210600, 828211500, 828212400, 828213300, 828214200,
    828215100, 828216000, 828216900, 828217800, 828218700, 828219600,
    828220500, 828221400, 828222300, 828223200, 828224100, 828225000,
    828225900, 828226800, 828227700, 828228600, 828229500, 828230400,
    828231300, 828232200, 828233100, 828234000, 828234900, 828235800,
    828236700, 828237600, 828238500, 828239400, 828240300, 828241200,
    828242100, 828243000, 828243900, 828244800, 828245700, 828246600,
    828247500, 828248400, 828249300, 828250200, 828251100, 828252000,
    828252900, 828253800, 828254700, 828255600, 828256500, 828257400,
    828258300, 828259200, 828260100, 828261000, 828261900, 828262800,
    828263700, 828264600, 828265500, 828266400, 828267300, 828268200,
    828269100, 828270000, 828270900, 828271800, 828272700, 828273600,
    828274500, 828275400, 828276300, 828277200, 828278100, 828279000,
    828279900, 828280800, 828281700, 828282600, 828283500, 828284400,
    828285300, 828286200, 828287100, 828288000, 828288900, 828289800,
    828290700, 828291600, 828292500, 828293400, 828294300, 828295200,
    828296100, 828297000, 828297900, 828298800, 828299700, 828300600,
    828301500, 828302400, 828303300, 828304200, 828305100, 828306000,
    828306900, 828307800, 828308700, 828309600, 828310500, 828311400,
    828312300, 828313200, 828314100, 828315000, 828315900, 828316800,
    828317700, 828318600, 828319500, 828320400, 828321300, 828322200,
    828323100, 828324000, 828324900, 828325800, 828326700, 828327600,
    828328500, 828329400, 828330300, 828331200, 828332100, 828333000,
    828333900, 828334800, 828335700, 828336600, 828337500, 828338400,
    828339300, 828340200, 828341100, 828342000, 828342900, 828343800,
    828344700, 828345600, 828346500, 828347400, 828348300, 828349200,
    828350100, 828351000, 828351900, 828352800, 828353700, 828354600,
    828355500, 828356400, 828357300, 828358200, 828359100, 828360000,
    828360900, 828361800, 828362700, 828363600, 828364500, 828365400,
    828366300, 828367200, 828368100, 828369000, 828369900, 828370800,
    828371700, 828372600, 828373500, 828374400, 828375300, 828376200,
    828377100, 828378000, 828378900, 828379800, 828380700, 828381600,
    828382500, 828383400, 828384300, 828385200, 828386100, 828387000,
    828387900, 828388800, 828389700, 828390600, 828391500, 828392400,
    828393300, 828394200, 828395100, 828396000, 828396900, 828397800,
    828398700, 828399600, 828400500, 828401400, 828402300, 828403200,
    828404100, 828405000, 828405900, 828406800, 828407700, 828408600,
    828409500, 828410400, 828411300, 828412200, 828413100, 828414000,
    828414900, 828415800, 828416700, 828417600, 828418500, 828419400,
    828420300, 828421200, 828422100, 828423000, 828423900, 828424800,
    828425700, 828426600, 828427500, 828428400, 828429300, 828430200,
    828431100, 828432000, 828432900, 828433800, 828434700, 828435600,
    828436500, 828437400, 828438300, 828439200, 828440100, 828441000,
    828441900, 828442800, 828443700, 828444600, 828445500, 828446400,
    828447300, 828448200, 828449100, 828450000, 828450900, 828451800,
    828452700, 828453600, 828454500, 828455400, 828456300, 828457200,
    828458100, 828459000, 828459900, 828460800, 828461700, 828462600,
    828463500, 828464400, 828465300, 828466200, 828467100, 828468000,
    828468900, 828469800, 828470700, 828471600, 828472500, 828473400,
    828474300, 828475200, 828476100, 828477000, 828477900, 828478800,
    828479700, 828480600, 828481500, 828482400, 828483300, 828484200,
    828485100, 828486000, 828486900, 828487800, 828488700, 828489600,
    828490500, 828491400, 828492300, 828493200, 828494100, 828495000,
    828495900, 828496800, 828497700, 828498600, 828499500, 828500400,
    828501300, 828502200, 828503100, 828504000, 828504900, 828505800,
    828506700, 828507600, 828508500, 828509400, 828510300, 828511200,
    828512100, 828513000, 828513900, 828514800, 828515700, 828516600,
    828517500, 828518400, 828519300, 828520200, 828521100, 828522000,
    828522900, 828523800, 828524700, 828525600, 828526500, 828527400,
    828528300, 828529200, 828530100, 828531000, 828531900, 828532800,
    828533700, 828534600, 828535500, 828536400, 828537300, 828538200,
    828539100, 828540000, 828540900, 828541800, 828542700, 828543600,
    828544500, 828545400, 828546300, 828547200, 828548100, 828549000,
    828549900, 828550800, 828551700, 828552600, 828553500, 828554400,
    828555300, 828556200, 828557100, 828558000, 828558900, 828559800,
    828560700, 828561600, 828562500, 828563400, 828564300, 828565200,
    828566100, 828567000, 828567900, 828568800, 828569700, 828570600,
    828571500, 828572400, 828573300, 828574200, 828575100, 828576000,
    828576900, 828577800, 828578700, 828579600, 828580500, 828581400,
    828582300, 828583200, 828584100, 828585000, 828585900, 828586800,
    828587700, 828588600, 828589500, 828590400, 828591300, 828592200,
    828593100, 828594000, 828594900, 828595800, 828596700, 828597600,
    828598500, 828599400, 828600300, 828601200, 828602100, 828603000,
    828603900, 828604800, 828605700, 828606600, 828607500, 828608400,
    828609300, 828610200, 828611100, 828612000, 828612900, 828613800,
    828614700, 828615600, 828616500, 828617400, 828618300, 828619200,
    828620100, 828621000, 828621900, 828622800, 828623700, 828624600,
    828625500, 828626400, 828627300, 828628200, 828629100, 828630000,
    828630900, 828631800, 828632700, 828633600, 828634500, 828635400,
    828636300, 828637200, 828638100, 828639000, 828639900, 828640800,
    828641700, 828642600, 828643500, 828644400, 828645300, 828646200,
    828647100, 828648000, 828648900, 828649800, 828650700, 828651600,
    828652500, 828653400, 828654300, 828655200, 828656100, 828657000,
    828657900, 828658800, 828659700, 828660600, 828661500, 828662400,
    828663300, 828664200, 828665100, 828666000, 828666900, 828667800,
    828668700, 828669600, 828670500, 828671400, 828672300, 828673200,
    828674100, 828675000, 828675900, 828676800, 828677700, 828678600,
    828679500, 828680400, 828681300, 828682200, 828683100, 828684000,
    828684900, 828685800, 828686700, 828687600, 828688500, 828689400,
    828690300, 828691200, 828692100, 828693000, 828693900, 828694800,
    828695700, 828696600, 828697500, 828698400, 828699300, 828700200,
    828701100, 828702000, 828702900, 828703800, 828704700, 828705600,
    828706500, 828707400, 828708300, 828709200, 828710100, 828711000,
    828711900, 828712800, 828713700, 828714600, 828715500, 828716400,
    828717300, 828718200, 828719100, 828720000, 828720900, 828721800,
    828722700, 828723600, 828724500, 828725400, 828726300, 828727200,
    828728100, 828729000, 828729900, 828730800, 828731700, 828732600,
    828733500, 828734400, 828735300, 828736200, 828737100, 828738000,
    828738900, 828739800, 828740700, 828741600, 828742500, 828743400,
    828744300, 828745200, 828746100, 828747000, 828747900, 828748800,
    828749700, 828750600, 828751500, 828752400, 828753300, 828754200,
    828755100, 828756000, 828756900, 828757800, 828758700, 828759600,
    828760500, 828761400, 828762300, 828763200, 828764100, 828765000,
    828765900, 828766800, 828767700, 828768600, 828769500, 828770400,
    828771300, 828772200, 828773100, 828774000, 828774900, 828775800,
    828776700, 828777600, 828778500, 828779400, 828780300, 828781200,
    828782100, 828783000, 828783900, 828784800, 828785700, 828786600,
    828787500, 828788400, 828789300, 828790200, 828791100, 828792000,
    828792900, 828793800, 828794700, 828795600, 828796500, 828797400,
    828798300, 828799200, 828800100, 828801000, 828801900, 828802800,
    828803700, 828804600, 828805500, 828806400, 828807300, 828808200,
    828809100, 828810000, 828810900, 828811800, 828812700, 828813600,
    828814500, 828815400, 828816300, 828817200, 828818100, 828819000,
    828819900, 828820800, 828821700, 828822600, 828823500, 828824400,
    828825300, 828826200, 828827100, 828828000, 828828900, 828829800,
    828830700, 828831600, 828832500, 828833400, 828834300, 828835200,
    828836100, 828837000, 828837900, 828838800, 828839700, 828840600,
    828841500, 828842400, 828843300, 828844200, 828845100, 828846000,
    828846900, 828847800, 828848700, 828849600, 828850500, 828851400,
    828852300, 828853200, 828854100, 828855000, 828855900, 828856800,
    828857700, 828858600, 828859500, 828860400, 828861300, 828862200,
    828863100, 828864000, 828864900, 828865800, 828866700, 828867600,
    828868500, 828869400, 828870300, 828871200, 828872100, 828873000,
    828873900, 828874800, 828875700, 828876600, 828877500, 828878400,
    828879300, 828880200, 828881100, 828882000, 828882900, 828883800,
    828884700, 828885600, 828886500, 828887400, 828888300, 828889200,
    828890100, 828891000, 828891900, 828892800, 828893700, 828894600,
    828895500, 828896400, 828897300, 828898200, 828899100, 828900000,
    828900900, 828901800, 828902700, 828903600, 828904500, 828905400,
    828906300, 828907200, 828908100, 828909000, 828909900, 828910800,
    828911700, 828912600, 828913500, 828914400, 828915300, 828916200,
    828917100, 828918000, 828918900, 828919800, 828920700, 828921600,
    828922500, 828923400, 828924300, 828925200, 828926100, 828927000,
    828927900, 828928800, 828929700, 828930600, 828931500, 828932400,
    828933300, 828934200, 828935100, 828936000, 828936900, 828937800,
    828938700, 828939600, 828940500, 828941400, 828942300, 828943200,
    828944100, 828945000, 828945900, 828946800, 828947700, 828948600,
    828949500, 828950400, 828951300, 828952200, 828953100, 828954000,
    828954900, 828955800, 828956700, 828957600, 828958500, 828959400,
    828960300, 828961200, 828962100, 828963000, 828963900, 828964800,
    828965700, 828966600, 828967500, 828968400, 828969300, 828970200,
    828971100, 828972000, 828972900, 828973800, 828974700, 828975600,
    828976500, 828977400, 828978300, 828979200, 828980100, 828981000,
    828981900, 828982800, 828983700, 828984600, 828985500, 828986400,
    828987300, 828988200, 828989100, 828990000, 828990900, 828991800,
    828992700, 828993600, 828994500, 828995400, 828996300, 828997200,
    828998100, 828999000, 828999900, 829000800, 829001700, 829002600,
    829003500, 829004400, 829005300, 829006200, 829007100, 829008000,
    829008900, 829009800, 829010700, 829011600, 829012500, 829013400,
    829014300, 829015200, 829016100, 829017000, 829017900, 829018800,
    829019700, 829020600, 829021500, 829022400, 829023300, 829024200,
    829025100, 829026000, 829026900, 829027800, 829028700, 829029600,
    829030500, 829031400, 829032300, 829033200, 829034100, 829035000,
    829035900, 829036800, 829037700, 829038600, 829039500, 829040400,
    829041300, 829042200, 829043100, 829044000, 829044900, 829045800,
    829046700, 829047600, 829048500, 829049400, 829050300, 829051200,
    829052100, 829053000, 829053900, 829054800, 829055700, 829056600,
    829057500, 829058400, 829059300, 829060200, 829061100, 829062000,
    829062900, 829063800, 829064700, 829065600, 829066500, 829067400,
    829068300, 829069200, 829070100, 829071000, 829071900, 829072800,
    829073700, 829074600, 829075500, 829076400, 829077300, 829078200,
    829079100, 829080000, 829080900, 829081800, 829082700, 829083600,
    829084500, 829085400, 829086300, 829087200, 829088100, 829089000,
    829089900, 829090800, 829091700, 829092600, 829093500, 829094400,
    829095300, 829096200, 829097100, 829098000, 829098900, 829099800,
    829100700, 829101600, 829102500, 829103400, 829104300, 829105200,
    829106100, 829107000, 829107900, 829108800, 829109700, 829110600,
    829111500, 829112400, 829113300, 829114200, 829115100, 829116000,
    829116900, 829117800, 829118700, 829119600, 829120500, 829121400,
    829122300, 829123200, 829124100, 829125000, 829125900, 829126800,
    829127700, 829128600, 829129500, 829130400, 829131300, 829132200,
    829133100, 829134000, 829134900, 829135800, 829136700, 829137600,
    829138500, 829139400, 829140300, 829141200, 829142100, 829143000,
    829143900, 829144800, 829145700, 829146600, 829147500, 829148400,
    829149300, 829150200, 829151100, 829152000, 829152900, 829153800,
    829154700, 829155600, 829156500, 829157400, 829158300, 829159200,
    829160100, 829161000, 829161900, 829162800, 829163700, 829164600,
    829165500, 829166400, 829167300, 829168200, 829169100, 829170000,
    829170900, 829171800, 829172700, 829173600, 829174500, 829175400,
    829176300, 829177200, 829178100, 829179000, 829179900, 829180800,
    829181700, 829182600, 829183500, 829184400, 829185300, 829186200,
    829187100, 829188000, 829188900, 829189800, 829190700, 829191600,
    829192500, 829193400, 829194300, 829195200, 829196100, 829197000,
    829197900, 829198800, 829199700, 829200600, 829201500, 829202400,
    829203300, 829204200, 829205100, 829206000, 829206900, 829207800,
    829208700, 829209600, 829210500, 829211400, 829212300, 829213200,
    829214100, 829215000, 829215900, 829216800, 829217700, 829218600,
    829219500, 829220400, 829221300, 829222200, 829223100, 829224000,
    829224900, 829225800, 829226700, 829227600, 829228500, 829229400,
    829230300, 829231200, 829232100, 829233000, 829233900, 829234800,
    829235700, 829236600, 829237500, 829238400, 829239300, 829240200,
    829241100, 829242000, 829242900, 829243800, 829244700, 829245600,
    829246500, 829247400, 829248300, 829249200, 829250100, 829251000,
    829251900, 829252800, 829253700, 829254600, 829255500, 829256400,
    829257300, 829258200, 829259100, 829260000, 829260900, 829261800,
    829262700, 829263600, 829264500, 829265400, 829266300, 829267200,
    829268100, 829269000, 829269900, 829270800, 829271700, 829272600,
    829273500, 829274400, 829275300, 829276200, 829277100, 829278000,
    829278900, 829279800, 829280700, 829281600, 829282500, 829283400,
    829284300, 829285200, 829286100, 829287000, 829287900, 829288800,
    829289700, 829290600, 829291500, 829292400, 829293300, 829294200,
    829295100, 829296000, 829296900, 829297800, 829298700, 829299600,
    829300500, 829301400, 829302300, 829303200, 829304100, 829305000,
    829305900, 829306800, 829307700, 829308600, 829309500, 829310400,
    829311300, 829312200, 829313100, 829314000, 829314900, 829315800,
    829316700, 829317600, 829318500, 829319400, 829320300, 829321200,
    829322100, 829323000, 829323900, 829324800, 829325700, 829326600,
    829327500, 829328400, 829329300, 829330200, 829331100, 829332000,
    829332900, 829333800, 829334700, 829335600, 829336500, 829337400,
    829338300, 829339200, 829340100, 829341000, 829341900, 829342800,
    829343700, 829344600, 829345500, 829346400, 829347300, 829348200,
    829349100, 829350000, 829350900, 829351800, 829352700, 829353600,
    829354500, 829355400, 829356300, 829357200, 829358100, 829359000,
    829359900, 829360800, 829361700, 829362600, 829363500, 829364400,
    829365300, 829366200, 829367100, 829368000, 829368900, 829369800,
    829370700, 829371600, 829372500, 829373400, 829374300, 829375200,
    829376100, 829377000, 829377900, 829378800, 829379700, 829380600,
    829381500, 829382400, 829383300, 829384200, 829385100, 829386000,
    829386900, 829387800, 829388700, 829389600, 829390500, 829391400,
    829392300, 829393200, 829394100, 829395000, 829395900, 829396800,
    829397700, 829398600, 829399500, 829400400, 829401300, 829402200,
    829403100, 829404000, 829404900, 829405800, 829406700, 829407600,
    829408500, 829409400, 829410300, 829411200, 829412100, 829413000,
    829413900, 829414800, 829415700, 829416600, 829417500, 829418400,
    829419300, 829420200, 829421100, 829422000, 829422900, 829423800,
    829424700, 829425600, 829426500, 829427400, 829428300, 829429200,
    829430100, 829431000, 829431900, 829432800, 829433700, 829434600,
    829435500, 829436400, 829437300, 829438200, 829439100, 829440000,
    829440900, 829441800, 829442700, 829443600, 829444500, 829445400,
    829446300, 829447200, 829448100, 829449000, 829449900, 829450800,
    829451700, 829452600, 829453500, 829454400, 829455300, 829456200,
    829457100, 829458000, 829458900, 829459800, 829460700, 829461600,
    829462500, 829463400, 829464300, 829465200, 829466100, 829467000,
    829467900, 829468800, 829469700, 829470600, 829471500, 829472400,
    829473300, 829474200, 829475100, 829476000, 829476900, 829477800,
    829478700, 829479600, 829480500, 829481400, 829482300, 829483200,
    829484100, 829485000, 829485900, 829486800, 829487700, 829488600,
    829489500, 829490400, 829491300, 829492200, 829493100, 829494000,
    829494900, 829495800, 829496700, 829497600, 829498500, 829499400,
    829500300, 829501200, 829502100, 829503000, 829503900, 829504800,
    829505700, 829506600, 829507500, 829508400, 829509300, 829510200,
    829511100, 829512000, 829512900, 829513800, 829514700, 829515600,
    829516500, 829517400, 829518300, 829519200, 829520100, 829521000,
    829521900, 829522800, 829523700, 829524600, 829525500, 829526400,
    829527300, 829528200, 829529100, 829530000, 829530900, 829531800,
    829532700, 829533600, 829534500, 829535400, 829536300, 829537200,
    829538100, 829539000, 829539900, 829540800, 829541700, 829542600,
    829543500, 829544400, 829545300, 829546200, 829547100, 829548000,
    829548900, 829549800, 829550700, 829551600, 829552500, 829553400,
    829554300, 829555200, 829556100, 829557000, 829557900, 829558800,
    829559700, 829560600, 829561500, 829562400, 829563300, 829564200,
    829565100, 829566000, 829566900, 829567800, 829568700, 829569600,
    829570500, 829571400, 829572300, 829573200, 829574100, 829575000,
    829575900, 829576800, 829577700, 829578600, 829579500, 829580400,
    829581300, 829582200, 829583100, 829584000, 829584900, 829585800,
    829586700, 829587600, 829588500, 829589400, 829590300, 829591200,
    829592100, 829593000, 829593900, 829594800, 829595700, 829596600,
    829597500, 829598400, 829599300, 829600200, 829601100, 829602000,
    829602900, 829603800, 829604700, 829605600, 829606500, 829607400,
    829608300, 829609200, 829610100, 829611000, 829611900, 829612800,
    829613700, 829614600, 829615500, 829616400, 829617300, 829618200,
    829619100, 829620000, 829620900, 829621800, 829622700, 829623600,
    829624500, 829625400, 829626300, 829627200, 829628100, 829629000,
    829629900, 829630800, 829631700, 829632600, 829633500, 829634400,
    829635300, 829636200, 829637100, 829638000, 829638900, 829639800,
    829640700, 829641600, 829642500, 829643400, 829644300, 829645200,
    829646100, 829647000, 829647900, 829648800, 829649700, 829650600,
    829651500, 829652400, 829653300, 829654200, 829655100, 829656000,
    829656900, 829657800, 829658700, 829659600, 829660500, 829661400,
    829662300, 829663200, 829664100, 829665000, 829665900, 829666800,
    829667700, 829668600, 829669500, 829670400, 829671300, 829672200,
    829673100, 829674000, 829674900, 829675800, 829676700, 829677600,
    829678500, 829679400, 829680300, 829681200, 829682100, 829683000,
    829683900, 829684800, 829685700, 829686600, 829687500, 829688400,
    829689300, 829690200, 829691100, 829692000, 829692900, 829693800,
    829694700, 829695600, 829696500, 829697400, 829698300, 829699200,
    829700100, 829701000, 829701900, 829702800, 829703700, 829704600,
    829705500, 829706400, 829707300, 829708200, 829709100, 829710000,
    829710900, 829711800, 829712700, 829713600, 829714500, 829715400,
    829716300, 829717200, 829718100, 829719000, 829719900, 829720800,
    829721700, 829722600, 829723500, 829724400, 829725300, 829726200,
    829727100, 829728000, 829728900, 829729800, 829730700, 829731600,
    829732500, 829733400, 829734300, 829735200, 829736100, 829737000,
    829737900, 829738800, 829739700, 829740600, 829741500, 829742400,
    829743300, 829744200, 829745100, 829746000, 829746900, 829747800,
    829748700, 829749600, 829750500, 829751400, 829752300, 829753200,
    829754100, 829755000, 829755900, 829756800, 829757700, 829758600,
    829759500, 829760400, 829761300, 829762200, 829763100, 829764000,
    829764900, 829765800, 829766700, 829767600, 829768500, 829769400,
    829770300, 829771200, 829772100, 829773000, 829773900, 829774800,
    829775700, 829776600, 829777500, 829778400, 829779300, 829780200,
    829781100, 829782000, 829782900, 829783800, 829784700, 829785600,
    829786500, 829787400, 829788300, 829789200, 829790100, 829791000,
    829791900, 829792800, 829793700, 829794600, 829795500, 829796400,
    829797300, 829798200, 829799100, 829800000, 829800900, 829801800,
    829802700, 829803600, 829804500, 829805400, 829806300, 829807200,
    829808100, 829809000, 829809900, 829810800, 829811700, 829812600,
    829813500, 829814400, 829815300, 829816200, 829817100, 829818000,
    829818900, 829819800, 829820700, 829821600, 829822500, 829823400,
    829824300, 829825200, 829826100, 829827000, 829827900, 829828800,
    829829700, 829830600, 829831500, 829832400, 829833300, 829834200,
    829835100, 829836000, 829836900, 829837800, 829838700, 829839600,
    829840500, 829841400, 829842300, 829843200, 829844100, 829845000,
    829845900, 829846800, 829847700, 829848600, 829849500, 829850400,
    829851300, 829852200, 829853100, 829854000, 829854900, 829855800,
    829856700, 829857600, 829858500, 829859400, 829860300, 829861200,
    829862100, 829863000, 829863900, 829864800, 829865700, 829866600,
    829867500, 829868400, 829869300, 829870200, 829871100, 829872000,
    829872900, 829873800, 829874700, 829875600, 829876500, 829877400,
    829878300, 829879200, 829880100, 829881000, 829881900, 829882800,
    829883700, 829884600, 829885500, 829886400, 829887300, 829888200,
    829889100, 829890000, 829890900, 829891800, 829892700, 829893600,
    829894500, 829895400, 829896300, 829897200, 829898100, 829899000,
    829899900, 829900800, 829901700, 829902600, 829903500, 829904400,
    829905300, 829906200, 829907100, 829908000, 829908900, 829909800,
    829910700, 829911600, 829912500, 829913400, 829914300, 829915200,
    829916100, 829917000, 829917900, 829918800, 829919700, 829920600,
    829921500, 829922400, 829923300, 829924200, 829925100, 829926000,
    829926900, 829927800, 829928700, 829929600, 829930500, 829931400,
    829932300, 829933200, 829934100, 829935000, 829935900, 829936800,
    829937700, 829938600, 829939500, 829940400, 829941300, 829942200,
    829943100, 829944000, 829944900, 829945800, 829946700, 829947600,
    829948500, 829949400, 829950300, 829951200, 829952100, 829953000,
    829953900, 829954800, 829955700, 829956600, 829957500, 829958400,
    829959300, 829960200, 829961100, 829962000, 829962900, 829963800,
    829964700, 829965600, 829966500, 829967400, 829968300, 829969200,
    829970100, 829971000, 829971900, 829972800, 829973700, 829974600,
    829975500, 829976400, 829977300, 829978200, 829979100, 829980000,
    829980900, 829981800, 829982700, 829983600, 829984500, 829985400,
    829986300, 829987200, 829988100, 829989000, 829989900, 829990800,
    829991700, 829992600, 829993500, 829994400, 829995300, 829996200,
    829997100, 829998000, 829998900, 829999800, 830000700, 830001600,
    830002500, 830003400, 830004300, 830005200, 830006100, 830007000,
    830007900, 830008800, 830009700, 830010600, 830011500, 830012400,
    830013300, 830014200, 830015100, 830016000, 830016900, 830017800,
    830018700, 830019600, 830020500, 830021400, 830022300, 830023200,
    830024100, 830025000, 830025900, 830026800, 830027700, 830028600,
    830029500, 830030400, 830031300, 830032200, 830033100, 830034000,
    830034900, 830035800, 830036700, 830037600, 830038500, 830039400,
    830040300, 830041200, 830042100, 830043000, 830043900, 830044800,
    830045700, 830046600, 830047500, 830048400, 830049300, 830050200,
    830051100, 830052000, 830052900, 830053800, 830054700, 830055600,
    830056500, 830057400, 830058300, 830059200, 830060100, 830061000,
    830061900, 830062800, 830063700, 830064600, 830065500, 830066400,
    830067300, 830068200, 830069100, 830070000, 830070900, 830071800,
    830072700, 830073600, 830074500, 830075400, 830076300, 830077200,
    830078100, 830079000, 830079900, 830080800, 830081700, 830082600,
    830083500, 830084400, 830085300, 830086200, 830087100, 830088000,
    830088900, 830089800, 830090700, 830091600, 830092500, 830093400,
    830094300, 830095200, 830096100, 830097000, 830097900, 830098800,
    830099700, 830100600, 830101500, 830102400, 830103300, 830104200,
    830105100, 830106000, 830106900, 830107800, 830108700, 830109600,
    830110500, 830111400, 830112300, 830113200, 830114100, 830115000,
    830115900, 830116800, 830117700, 830118600, 830119500, 830120400,
    830121300, 830122200, 830123100, 830124000, 830124900, 830125800,
    830126700, 830127600, 830128500, 830129400, 830130300, 830131200,
    830132100, 830133000, 830133900, 830134800, 830135700, 830136600,
    830137500, 830138400, 830139300, 830140200, 830141100, 830142000,
    830142900, 830143800, 830144700, 830145600, 830146500, 830147400,
    830148300, 830149200, 830150100, 830151000, 830151900, 830152800,
    830153700, 830154600, 830155500, 830156400, 830157300, 830158200,
    830159100, 830160000, 830160900, 830161800, 830162700, 830163600,
    830164500, 830165400, 830166300, 830167200, 830168100, 830169000,
    830169900, 830170800, 830171700, 830172600, 830173500, 830174400,
    830175300, 830176200, 830177100, 830178000, 830178900, 830179800,
    830180700, 830181600, 830182500, 830183400, 830184300, 830185200,
    830186100, 830187000, 830187900, 830188800, 830189700, 830190600,
    830191500, 830192400, 830193300, 830194200, 830195100, 830196000,
    830196900, 830197800, 830198700, 830199600, 830200500, 830201400,
    830202300, 830203200, 830204100, 830205000, 830205900, 830206800,
    830207700, 830208600, 830209500, 830210400, 830211300, 830212200,
    830213100, 830214000, 830214900, 830215800, 830216700, 830217600,
    830218500, 830219400, 830220300, 830221200, 830222100, 830223000,
    830223900, 830224800, 830225700, 830226600, 830227500, 830228400,
    830229300, 830230200, 830231100, 830232000, 830232900, 830233800,
    830234700, 830235600, 830236500, 830237400, 830238300, 830239200,
    830240100, 830241000, 830241900, 830242800, 830243700, 830244600,
    830245500, 830246400, 830247300, 830248200, 830249100, 830250000,
    830250900, 830251800, 830252700, 830253600, 830254500, 830255400,
    830256300, 830257200, 830258100, 830259000, 830259900, 830260800,
    830261700, 830262600, 830263500, 830264400, 830265300, 830266200,
    830267100, 830268000, 830268900, 830269800, 830270700, 830271600,
    830272500, 830273400, 830274300, 830275200, 830276100, 830277000,
    830277900, 830278800, 830279700, 830280600, 830281500, 830282400,
    830283300, 830284200, 830285100, 830286000, 830286900, 830287800,
    830288700, 830289600, 830290500, 830291400, 830292300, 830293200,
    830294100, 830295000, 830295900, 830296800, 830297700, 830298600,
    830299500, 830300400, 830301300, 830302200, 830303100, 830304000,
    830304900, 830305800, 830306700, 830307600, 830308500, 830309400,
    830310300, 830311200, 830312100, 830313000, 830313900, 830314800,
    830315700, 830316600, 830317500, 830318400, 830319300, 830320200,
    830321100, 830322000, 830322900, 830323800, 830324700, 830325600,
    830326500, 830327400, 830328300, 830329200, 830330100, 830331000,
    830331900, 830332800, 830333700, 830334600, 830335500, 830336400,
    830337300, 830338200, 830339100, 830340000, 830340900, 830341800,
    830342700, 830343600, 830344500, 830345400, 830346300, 830347200,
    830348100, 830349000, 830349900, 830350800, 830351700, 830352600,
    830353500, 830354400, 830355300, 830356200, 830357100, 830358000,
    830358900, 830359800, 830360700, 830361600, 830362500, 830363400,
    830364300, 830365200, 830366100, 830367000, 830367900, 830368800,
    830369700, 830370600, 830371500, 830372400, 830373300, 830374200,
    830375100, 830376000, 830376900, 830377800, 830378700, 830379600,
    830380500, 830381400, 830382300, 830383200, 830384100, 830385000,
    830385900, 830386800, 830387700, 830388600, 830389500, 830390400,
    830391300, 830392200, 830393100, 830394000, 830394900, 830395800,
    830396700, 830397600, 830398500, 830399400, 830400300, 830401200,
    830402100, 830403000, 830403900, 830404800, 830405700, 830406600,
    830407500, 830408400, 830409300, 830410200, 830411100, 830412000,
    830412900, 830413800, 830414700, 830415600, 830416500, 830417400,
    830418300, 830419200, 830420100, 830421000, 830421900, 830422800,
    830423700, 830424600, 830425500, 830426400, 830427300, 830428200,
    830429100, 830430000, 830430900, 830431800, 830432700, 830433600,
    830434500, 830435400, 830436300, 830437200, 830438100, 830439000,
    830439900, 830440800, 830441700, 830442600, 830443500, 830444400,
    830445300, 830446200, 830447100, 830448000, 830448900, 830449800,
    830450700, 830451600, 830452500, 830453400, 830454300, 830455200,
    830456100, 830457000, 830457900, 830458800, 830459700, 830460600,
    830461500, 830462400, 830463300, 830464200, 830465100, 830466000,
    830466900, 830467800, 830468700, 830469600, 830470500, 830471400,
    830472300, 830473200, 830474100, 830475000, 830475900, 830476800,
    830477700, 830478600, 830479500, 830480400, 830481300, 830482200,
    830483100, 830484000, 830484900, 830485800, 830486700, 830487600,
    830488500, 830489400, 830490300, 830491200, 830492100, 830493000,
    830493900, 830494800, 830495700, 830496600, 830497500, 830498400,
    830499300, 830500200, 830501100, 830502000, 830502900, 830503800,
    830504700, 830505600, 830506500, 830507400, 830508300, 830509200,
    830510100, 830511000, 830511900, 830512800, 830513700, 830514600,
    830515500, 830516400, 830517300, 830518200, 830519100, 830520000,
    830520900, 830521800, 830522700, 830523600, 830524500, 830525400,
    830526300, 830527200, 830528100, 830529000, 830529900, 830530800,
    830531700, 830532600, 830533500, 830534400, 830535300, 830536200,
    830537100, 830538000, 830538900, 830539800, 830540700, 830541600,
    830542500, 830543400, 830544300, 830545200, 830546100, 830547000,
    830547900, 830548800, 830549700, 830550600, 830551500, 830552400,
    830553300, 830554200, 830555100, 830556000, 830556900, 830557800,
    830558700, 830559600, 830560500, 830561400, 830562300, 830563200,
    830564100, 830565000, 830565900, 830566800, 830567700, 830568600,
    830569500, 830570400, 830571300, 830572200, 830573100, 830574000,
    830574900, 830575800, 830576700, 830577600, 830578500, 830579400,
    830580300, 830581200, 830582100, 830583000, 830583900, 830584800,
    830585700, 830586600, 830587500, 830588400, 830589300, 830590200,
    830591100, 830592000, 830592900, 830593800, 830594700, 830595600,
    830596500, 830597400, 830598300, 830599200, 830600100, 830601000,
    830601900, 830602800, 830603700, 830604600, 830605500, 830606400,
    830607300, 830608200, 830609100, 830610000, 830610900, 830611800,
    830612700, 830613600, 830614500, 830615400, 830616300, 830617200,
    830618100, 830619000, 830619900, 830620800, 830621700, 830622600,
    830623500, 830624400, 830625300, 830626200, 830627100, 830628000,
    830628900, 830629800, 830630700, 830631600, 830632500, 830633400,
    830634300, 830635200, 830636100, 830637000, 830637900, 830638800,
    830639700, 830640600, 830641500, 830642400, 830643300, 830644200,
    830645100, 830646000, 830646900, 830647800, 830648700, 830649600,
    830650500, 830651400, 830652300, 830653200, 830654100, 830655000,
    830655900, 830656800, 830657700, 830658600, 830659500, 830660400,
    830661300, 830662200, 830663100, 830664000, 830664900, 830665800,
    830666700, 830667600, 830668500, 830669400, 830670300, 830671200,
    830672100, 830673000, 830673900, 830674800, 830675700, 830676600,
    830677500, 830678400, 830679300, 830680200, 830681100, 830682000,
    830682900, 830683800, 830684700, 830685600, 830686500, 830687400,
    830688300, 830689200, 830690100, 830691000, 830691900, 830692800,
    830693700, 830694600, 830695500, 830696400, 830697300, 830698200,
    830699100, 830700000, 830700900, 830701800, 830702700, 830703600,
    830704500, 830705400, 830706300, 830707200, 830708100, 830709000,
    830709900, 830710800, 830711700, 830712600, 830713500, 830714400,
    830715300, 830716200, 830717100, 830718000, 830718900, 830719800,
    830720700, 830721600, 830722500, 830723400, 830724300, 830725200,
    830726100, 830727000, 830727900, 830728800, 830729700, 830730600,
    830731500, 830732400, 830733300, 830734200, 830735100, 830736000,
    830736900, 830737800, 830738700, 830739600, 830740500, 830741400,
    830742300, 830743200, 830744100, 830745000, 830745900, 830746800,
    830747700, 830748600, 830749500, 830750400, 830751300, 830752200,
    830753100, 830754000, 830754900, 830755800, 830756700, 830757600,
    830758500, 830759400, 830760300, 830761200, 830762100, 830763000,
    830763900, 830764800, 830765700, 830766600, 830767500, 830768400,
    830769300, 830770200, 830771100, 830772000, 830772900, 830773800,
    830774700, 830775600, 830776500, 830777400, 830778300, 830779200,
    830780100, 830781000, 830781900, 830782800, 830783700, 830784600,
    830785500, 830786400, 830787300, 830788200, 830789100, 830790000,
    830790900, 830791800, 830792700, 830793600, 830794500, 830795400,
    830796300, 830797200, 830798100, 830799000, 830799900, 830800800,
    830801700, 830802600, 830803500, 830804400, 830805300, 830806200,
    830807100, 830808000, 830808900, 830809800, 830810700, 830811600,
    830812500, 830813400, 830814300, 830815200, 830816100, 830817000,
    830817900, 830818800, 830819700, 830820600, 830821500, 830822400,
    830823300, 830824200, 830825100, 830826000, 830826900, 830827800,
    830828700, 830829600, 830830500, 830831400, 830832300, 830833200,
    830834100, 830835000, 830835900, 830836800, 830837700, 830838600,
    830839500, 830840400, 830841300, 830842200, 830843100, 830844000,
    830844900, 830845800, 830846700, 830847600, 830848500, 830849400,
    830850300, 830851200, 830852100, 830853000, 830853900, 830854800,
    830855700, 830856600, 830857500, 830858400, 830859300, 830860200,
    830861100, 830862000, 830862900, 830863800, 830864700, 830865600,
    830866500, 830867400, 830868300, 830869200, 830870100, 830871000,
    830871900, 830872800, 830873700, 830874600, 830875500, 830876400,
    830877300, 830878200, 830879100, 830880000, 830880900, 830881800,
    830882700, 830883600, 830884500, 830885400, 830886300, 830887200,
    830888100, 830889000, 830889900, 830890800, 830891700, 830892600,
    830893500, 830894400, 830895300, 830896200, 830897100, 830898000,
    830898900, 830899800, 830900700, 830901600, 830902500, 830903400,
    830904300, 830905200, 830906100, 830907000, 830907900, 830908800,
    830909700, 830910600, 830911500, 830912400, 830913300, 830914200,
    830915100, 830916000, 830916900, 830917800, 830918700, 830919600,
    830920500, 830921400, 830922300, 830923200, 830924100, 830925000,
    830925900, 830926800, 830927700, 830928600, 830929500, 830930400,
    830931300, 830932200, 830933100, 830934000, 830934900, 830935800,
    830936700, 830937600, 830938500, 830939400, 830940300, 830941200,
    830942100, 830943000, 830943900, 830944800, 830945700, 830946600,
    830947500, 830948400, 830949300, 830950200, 830951100, 830952000,
    830952900, 830953800, 830954700, 830955600, 830956500, 830957400,
    830958300, 830959200, 830960100, 830961000, 830961900, 830962800,
    830963700, 830964600, 830965500, 830966400, 830967300, 830968200,
    830969100, 830970000, 830970900, 830971800, 830972700, 830973600,
    830974500, 830975400, 830976300, 830977200, 830978100, 830979000,
    830979900, 830980800, 830981700, 830982600, 830983500, 830984400,
    830985300, 830986200, 830987100, 830988000, 830988900, 830989800,
    830990700, 830991600, 830992500, 830993400, 830994300, 830995200,
    830996100, 830997000, 830997900, 830998800, 830999700, 831000600,
    831001500, 831002400, 831003300, 831004200, 831005100, 831006000,
    831006900, 831007800, 831008700, 831009600, 831010500, 831011400,
    831012300, 831013200, 831014100, 831015000, 831015900, 831016800,
    831017700, 831018600, 831019500, 831020400, 831021300, 831022200,
    831023100, 831024000, 831024900, 831025800, 831026700, 831027600,
    831028500, 831029400, 831030300, 831031200, 831032100, 831033000,
    831033900, 831034800, 831035700, 831036600, 831037500, 831038400,
    831039300, 831040200, 831041100, 831042000, 831042900, 831043800,
    831044700, 831045600, 831046500, 831047400, 831048300, 831049200,
    831050100, 831051000, 831051900, 831052800, 831053700, 831054600,
    831055500, 831056400, 831057300, 831058200, 831059100, 831060000,
    831060900, 831061800, 831062700, 831063600, 831064500, 831065400,
    831066300, 831067200, 831068100, 831069000, 831069900, 831070800,
    831071700, 831072600, 831073500, 831074400, 831075300, 831076200,
    831077100, 831078000, 831078900, 831079800, 831080700, 831081600,
    831082500, 831083400, 831084300, 831085200, 831086100, 831087000,
    831087900, 831088800, 831089700, 831090600, 831091500, 831092400,
    831093300, 831094200, 831095100, 831096000, 831096900, 831097800,
    831098700, 831099600, 831100500, 831101400, 831102300, 831103200,
    831104100, 831105000, 831105900, 831106800, 831107700, 831108600,
    831109500, 831110400, 831111300, 831112200, 831113100, 831114000,
    831114900, 831115800, 831116700, 831117600, 831118500, 831119400,
    831120300, 831121200, 831122100, 831123000, 831123900, 831124800,
    831125700, 831126600, 831127500, 831128400, 831129300, 831130200,
    831131100, 831132000, 831132900, 831133800, 831134700, 831135600,
    831136500, 831137400, 831138300, 831139200, 831140100, 831141000,
    831141900, 831142800, 831143700, 831144600, 831145500, 831146400,
    831147300, 831148200, 831149100, 831150000, 831150900, 831151800,
    831152700, 831153600, 831154500, 831155400, 831156300, 831157200,
    831158100, 831159000, 831159900, 831160800, 831161700, 831162600,
    831163500, 831164400, 831165300, 831166200, 831167100, 831168000,
    831168900, 831169800, 831170700, 831171600, 831172500, 831173400,
    831174300, 831175200, 831176100, 831177000, 831177900, 831178800,
    831179700, 831180600, 831181500, 831182400, 831183300, 831184200,
    831185100, 831186000, 831186900, 831187800, 831188700, 831189600,
    831190500, 831191400, 831192300, 831193200, 831194100, 831195000,
    831195900, 831196800, 831197700, 831198600, 831199500, 831200400,
    831201300, 831202200, 831203100, 831204000, 831204900, 831205800,
    831206700, 831207600, 831208500, 831209400, 831210300, 831211200,
    831212100, 831213000, 831213900, 831214800, 831215700, 831216600,
    831217500, 831218400, 831219300, 831220200, 831221100, 831222000,
    831222900, 831223800, 831224700, 831225600, 831226500, 831227400,
    831228300, 831229200, 831230100, 831231000, 831231900, 831232800,
    831233700, 831234600, 831235500, 831236400, 831237300, 831238200,
    831239100, 831240000, 831240900, 831241800, 831242700, 831243600,
    831244500, 831245400, 831246300, 831247200, 831248100, 831249000,
    831249900, 831250800, 831251700, 831252600, 831253500, 831254400,
    831255300, 831256200, 831257100, 831258000, 831258900, 831259800,
    831260700, 831261600, 831262500, 831263400, 831264300, 831265200,
    831266100, 831267000, 831267900, 831268800, 831269700, 831270600,
    831271500, 831272400, 831273300, 831274200, 831275100, 831276000,
    831276900, 831277800, 831278700, 831279600, 831280500, 831281400,
    831282300, 831283200, 831284100, 831285000, 831285900, 831286800,
    831287700, 831288600, 831289500, 831290400, 831291300, 831292200,
    831293100, 831294000, 831294900, 831295800, 831296700, 831297600,
    831298500, 831299400, 831300300, 831301200, 831302100, 831303000,
    831303900, 831304800, 831305700, 831306600, 831307500, 831308400,
    831309300, 831310200, 831311100, 831312000, 831312900, 831313800,
    831314700, 831315600, 831316500, 831317400, 831318300, 831322800,
    831323700, 831324600, 831325500, 831326400, 831327300, 831328200,
    831329100, 831330000, 831330900, 831331800, 831332700, 831333600,
    831334500, 831335400, 831336300, 831337200, 831338100, 831339000,
    831339900, 831340800, 831341700, 831342600, 831343500, 831344400,
    831345300, 831346200, 831347100, 831348000, 831348900, 831349800,
    831350700, 831351600, 831352500, 831353400, 831354300, 831355200,
    831356100, 831357000, 831357900, 831358800, 831359700, 831360600,
    831361500, 831362400, 831363300, 831364200, 831365100, 831366000,
    831366900, 831367800, 831368700, 831369600, 831370500, 831371400,
    831372300, 831373200, 831374100, 831375000, 831375900, 831376800,
    831377700, 831378600, 831379500, 831380400, 831381300, 831382200,
    831383100, 831384000, 831384900, 831385800, 831386700, 831387600,
    831388500, 831389400, 831390300, 831391200, 831392100, 831393000,
    831393900, 831394800, 831395700, 831396600, 831397500, 831398400,
    831399300, 831400200, 831401100, 831402000, 831402900, 831403800,
    831404700, 831405600, 831406500, 831407400, 831408300, 831409200,
    831410100, 831411000, 831411900, 831412800, 831413700, 831414600,
    831415500, 831416400, 831417300, 831418200, 831419100, 831420000,
    831420900, 831421800, 831422700, 831423600, 831424500, 831425400,
    831426300, 831427200, 831428100, 831429000, 831429900, 831430800,
    831431700, 831432600, 831433500, 831434400, 831435300, 831436200,
    831437100, 831438000, 831438900, 831439800, 831440700, 831441600,
    831442500, 831443400, 831444300, 831445200, 831446100, 831447000,
    831447900, 831448800, 831449700, 831450600, 831451500, 831452400,
    831453300, 831454200, 831455100, 831456000, 831456900, 831457800,
    831458700, 831459600, 831460500, 831461400, 831462300, 831463200,
    831464100, 831465000, 831465900, 831466800, 831467700, 831468600,
    831469500, 831470400, 831471300, 831472200, 831473100, 831474000,
    831474900, 831475800, 831476700, 831477600, 831478500, 831479400,
    831480300, 831481200, 831482100, 831483000, 831483900, 831484800,
    831485700, 831486600, 831487500, 831488400, 831489300, 831490200,
    831491100, 831492000, 831492900, 831493800, 831494700, 831495600,
    831496500, 831497400, 831498300, 831499200, 831500100, 831501000,
    831501900, 831502800, 831503700, 831504600, 831505500, 831506400,
    831507300, 831508200, 831509100, 831510000, 831510900, 831511800,
    831512700, 831513600, 831514500, 831515400, 831516300, 831517200,
    831518100, 831519000, 831519900, 831520800, 831521700, 831522600,
    831523500, 831524400, 831525300, 831526200, 831527100, 831528000,
    831528900, 831529800, 831530700, 831531600, 831532500, 831533400,
    831534300, 831535200, 831536100, 831537000, 831537900, 831538800,
    831539700, 831540600, 831541500, 831542400, 831543300, 831544200,
    831545100, 831546000, 831546900, 831547800, 831548700, 831549600,
    831550500, 831551400, 831552300, 831553200, 831554100, 831555000,
    831555900, 831556800, 831557700, 831558600, 831559500, 831560400,
    831561300, 831562200, 831563100, 831564000, 831564900, 831565800,
    831566700, 831567600, 831568500, 831569400, 831570300, 831571200,
    831572100, 831573000, 831573900, 831574800, 831575700, 831576600,
    831577500, 831578400, 831579300, 831580200, 831581100, 831582000,
    831582900, 831583800, 831584700, 831585600, 831586500, 831587400,
    831588300, 831589200, 831590100, 831591000, 831591900, 831592800,
    831593700, 831594600, 831595500, 831596400, 831597300, 831598200,
    831599100, 831600000, 831600900, 831601800, 831602700, 831603600,
    831604500, 831605400, 831606300, 831607200, 831608100, 831609000,
    831609900, 831610800, 831611700, 831612600, 831613500, 831614400,
    831615300, 831616200, 831617100, 831618000, 831618900, 831619800,
    831620700, 831621600, 831622500, 831623400, 831624300, 831625200,
    831626100, 831627000, 831627900, 831628800, 831629700, 831630600,
    831631500, 831632400, 831633300, 831634200, 831635100, 831636000,
    831636900, 831637800, 831638700, 831639600, 831640500, 831641400,
    831642300, 831643200, 831644100, 831645000, 831645900, 831646800,
    831647700, 831648600, 831649500, 831650400, 831651300, 831652200,
    831653100, 831654000, 831654900, 831655800, 831656700, 831657600,
    831658500, 831659400, 831660300, 831661200, 831662100, 831663000,
    831663900, 831664800, 831665700, 831666600, 831667500, 831668400,
    831669300, 831670200, 831671100, 831672000, 831672900, 831673800,
    831674700, 831675600, 831676500, 831677400, 831678300, 831679200,
    831680100, 831681000, 831681900, 831682800, 831683700, 831684600,
    831685500, 831686400, 831687300, 831688200, 831689100, 831690000,
    831690900, 831691800, 831692700, 831693600, 831694500, 831695400,
    831696300, 831697200, 831698100, 831699000, 831699900, 831700800,
    831701700, 831702600, 831703500, 831704400, 831705300, 831706200,
    831707100, 831708000, 831708900, 831709800, 831710700, 831711600,
    831712500, 831713400, 831714300, 831715200, 831716100, 831717000,
    831717900, 831718800, 831719700, 831720600, 831721500, 831722400,
    831723300, 831724200, 831725100, 831726000, 831726900, 831727800,
    831728700, 831729600, 831730500, 831731400, 831732300, 831733200,
    831734100, 831735000, 831735900, 831736800, 831737700, 831738600,
    831739500, 831740400, 831741300, 831742200, 831743100, 831744000,
    831744900, 831745800, 831746700, 831747600, 831748500, 831749400,
    831750300, 831751200, 831752100, 831753000, 831753900, 831754800,
    831755700, 831756600, 831757500, 831758400, 831759300, 831760200,
    831761100, 831762000, 831762900, 831763800, 831764700, 831765600,
    831766500, 831767400, 831768300, 831769200, 831770100, 831771000,
    831771900, 831772800, 831773700, 831774600, 831775500, 831776400,
    831777300, 831778200, 831779100, 831780000, 831780900, 831781800,
    831782700, 831783600, 831784500, 831785400, 831786300, 831787200,
    831788100, 831789000, 831789900, 831790800, 831791700, 831792600,
    831793500, 831794400, 831795300, 831796200, 831797100, 831798000,
    831798900, 831799800, 831800700, 831801600, 831802500, 831803400,
    831804300, 831805200, 831806100, 831807000, 831807900, 831808800,
    831809700, 831810600, 831811500, 831812400, 831813300, 831814200,
    831815100, 831816000, 831816900, 831817800, 831818700, 831819600,
    831820500, 831821400, 831822300, 831823200, 831824100, 831825000,
    831825900, 831826800, 831827700, 831828600, 831829500, 831830400,
    831831300, 831832200, 831833100, 831834000, 831834900, 831835800,
    831836700, 831837600, 831838500, 831839400, 831840300, 831841200,
    831842100, 831843000, 831843900, 831844800, 831845700, 831846600,
    831847500, 831848400, 831849300, 831850200, 831851100, 831852000,
    831852900, 831853800, 831854700, 831855600, 831856500, 831857400,
    831858300, 831859200, 831860100, 831861000, 831861900, 831862800,
    831863700, 831864600, 831865500, 831866400, 831867300, 831868200,
    831869100, 831870000, 831870900, 831871800, 831872700, 831873600,
    831874500, 831875400, 831876300, 831877200, 831878100, 831879000,
    831879900, 831880800, 831881700, 831882600, 831883500, 831884400,
    831885300, 831886200, 831887100, 831888000, 831888900, 831889800,
    831890700, 831891600, 831892500, 831893400, 831894300, 831895200,
    831896100, 831897000, 831897900, 831898800, 831899700, 831900600,
    831901500, 831902400, 831903300, 831904200, 831905100, 831906000,
    831906900, 831907800, 831908700, 831909600, 831910500, 831911400,
    831912300, 831913200, 831914100, 831915000, 831915900, 831916800,
    831917700, 831918600, 831919500, 831920400, 831921300, 831922200,
    831923100, 831924000, 831924900, 831925800, 831926700, 831927600,
    831928500, 831929400, 831930300, 831931200, 831932100, 831933000,
    831933900, 831934800, 831935700, 831936600, 831937500, 831938400,
    831939300, 831940200, 831941100, 831942000, 831942900, 831943800,
    831944700, 831945600, 831946500, 831947400, 831948300, 831949200,
    831950100, 831951000, 831951900, 831952800, 831953700, 831954600,
    831955500, 831956400, 831957300, 831958200, 831959100, 831960000,
    831960900, 831961800, 831962700, 831963600, 831964500, 831965400,
    831966300, 831967200, 831968100, 831969000, 831969900, 831970800,
    831971700, 831972600, 831973500, 831974400, 831975300, 831976200,
    831977100, 831978000, 831978900, 831979800, 831980700, 831981600,
    831982500, 831983400, 831984300, 831985200, 831986100, 831987000,
    831987900, 831988800, 831989700, 831990600, 831991500, 831992400,
    831993300, 831994200, 831995100, 831996000, 831996900, 831997800,
    831998700, 831999600, 832000500, 832001400, 832002300, 832003200,
    832004100, 832005000, 832005900, 832006800, 832007700, 832008600,
    832009500, 832010400, 832011300, 832012200, 832013100, 832014000,
    832014900, 832015800, 832016700, 832017600, 832018500, 832019400,
    832020300, 832021200, 832022100, 832023000, 832023900, 832024800,
    832025700, 832026600, 832027500, 832028400, 832029300, 832030200,
    832031100, 832032000, 832032900, 832033800, 832034700, 832035600,
    832036500, 832037400, 832038300, 832039200, 832040100, 832041000,
    832041900, 832042800, 832043700, 832044600, 832045500, 832046400,
    832047300, 832048200, 832049100, 832050000, 832050900, 832051800,
    832052700, 832053600, 832054500, 832055400, 832056300, 832057200,
    832058100, 832059000, 832059900, 832060800, 832061700, 832062600,
    832063500, 832064400, 832065300, 832066200, 832067100, 832068000,
    832068900, 832069800, 832070700, 832071600, 832072500, 832073400,
    832074300, 832075200, 832076100, 832077000, 832077900, 832078800,
    832079700, 832080600, 832081500, 832082400, 832083300, 832084200,
    832085100, 832086000, 832086900, 832087800, 832088700, 832089600,
    832090500, 832091400, 832092300, 832093200, 832094100, 832095000,
    832095900, 832096800, 832097700, 832098600, 832099500, 832100400,
    832101300, 832102200, 832103100, 832104000, 832104900, 832105800,
    832106700, 832107600, 832108500, 832109400, 832110300, 832111200,
    832112100, 832113000, 832113900, 832114800, 832115700, 832116600,
    832117500, 832118400, 832119300, 832120200, 832121100, 832122000,
    832122900, 832123800, 832124700, 832125600, 832126500, 832127400,
    832128300, 832129200, 832130100, 832131000, 832131900, 832132800,
    832133700, 832134600, 832135500, 832136400, 832137300, 832138200,
    832139100, 832140000, 832140900, 832141800, 832142700, 832143600,
    832144500, 832145400, 832146300, 832147200, 832148100, 832149000,
    832149900, 832150800, 832151700, 832152600, 832153500, 832154400,
    832155300, 832156200, 832157100, 832158000, 832158900, 832159800,
    832160700, 832161600, 832162500, 832163400, 832164300, 832165200,
    832166100, 832167000, 832167900, 832168800, 832169700, 832170600,
    832171500, 832172400, 832173300, 832174200, 832175100, 832176000,
    832176900, 832177800, 832178700, 832179600, 832180500, 832181400,
    832182300, 832183200, 832184100, 832185000, 832185900, 832186800,
    832187700, 832188600, 832189500, 832190400, 832191300, 832192200,
    832193100, 832194000, 832194900, 832195800, 832196700, 832197600,
    832198500, 832199400, 832200300, 832201200, 832202100, 832203000,
    832203900, 832204800, 832205700, 832206600, 832207500, 832208400,
    832209300, 832210200, 832211100, 832212000, 832212900, 832213800,
    832214700, 832215600, 832216500, 832217400, 832218300, 832219200,
    832220100, 832221000, 832221900, 832222800, 832223700, 832224600,
    832225500, 832226400, 832227300, 832228200, 832229100, 832230000,
    832230900, 832231800, 832232700, 832233600, 832234500, 832235400,
    832236300, 832237200, 832238100, 832239000, 832239900, 832240800,
    832241700, 832242600, 832243500, 832244400, 832245300, 832246200,
    832247100, 832248000, 832248900, 832249800, 832250700, 832251600,
    832252500, 832253400, 832254300, 832255200, 832256100, 832257000,
    832257900, 832258800, 832259700, 832260600, 832261500, 832262400,
    832263300, 832264200, 832265100, 832266000, 832266900, 832267800,
    832268700, 832269600, 832270500, 832271400, 832272300, 832273200,
    832274100, 832275000, 832275900, 832276800, 832277700, 832278600,
    832279500, 832280400, 832281300, 832282200, 832283100, 832284000,
    832284900, 832285800, 832286700, 832287600, 832288500, 832289400,
    832290300, 832291200, 832292100, 832293000, 832293900, 832294800,
    832295700, 832296600, 832297500, 832298400, 832299300, 832300200,
    832301100, 832302000, 832302900, 832303800, 832304700, 832305600,
    832306500, 832307400, 832308300, 832309200, 832310100, 832311000,
    832311900, 832312800, 832313700, 832314600, 832315500, 832316400,
    832317300, 832318200, 832319100, 832320000, 832320900, 832321800,
    832322700, 832323600, 832324500, 832325400, 832326300, 832327200,
    832328100, 832329000, 832329900, 832330800, 832331700, 832332600,
    832333500, 832334400, 832335300, 832336200, 832337100, 832338000,
    832338900, 832339800, 832340700, 832341600, 832342500, 832343400,
    832344300, 832345200, 832346100, 832347000, 832347900, 832348800,
    832349700, 832350600, 832351500, 832352400, 832353300, 832354200,
    832355100, 832356000, 832356900, 832357800, 832358700, 832359600,
    832360500, 832361400, 832362300, 832363200, 832364100, 832365000,
    832365900, 832366800, 832367700, 832368600, 832369500, 832370400,
    832371300, 832372200, 832373100, 832374000, 832374900, 832375800,
    832376700, 832377600, 832378500, 832379400, 832380300, 832381200,
    832382100, 832383000, 832383900, 832384800, 832385700, 832386600,
    832387500, 832388400, 832389300, 832390200, 832391100, 832392000,
    832392900, 832393800, 832394700, 832395600, 832396500, 832397400,
    832398300, 832399200, 832400100, 832401000, 832401900, 832402800,
    832403700, 832404600, 832405500, 832406400, 832407300, 832408200,
    832409100, 832410000, 832410900, 832411800, 832412700, 832413600,
    832414500, 832415400, 832416300, 832417200, 832418100, 832419000,
    832419900, 832420800, 832421700, 832422600, 832423500, 832424400,
    832425300, 832426200, 832427100, 832428000, 832428900, 832429800,
    832430700, 832431600, 832432500, 832433400, 832434300, 832435200,
    832436100, 832437000, 832437900, 832438800, 832439700, 832440600,
    832441500, 832442400, 832443300, 832444200, 832445100, 832446000,
    832446900, 832447800, 832448700, 832449600, 832450500, 832451400,
    832452300, 832453200, 832454100, 832455000, 832455900, 832456800,
    832457700, 832458600, 832459500, 832460400, 832461300, 832462200,
    832463100, 832464000, 832464900, 832465800, 832466700, 832467600,
    832468500, 832469400, 832470300, 832471200, 832472100, 832473000,
    832473900, 832474800, 832475700, 832476600, 832477500, 832478400,
    832479300, 832480200, 832481100, 832482000, 832482900, 832483800,
    832484700, 832485600, 832486500, 832487400, 832488300, 832489200,
    832490100, 832491000, 832491900, 832492800, 832493700, 832494600,
    832495500, 832496400, 832497300, 832498200, 832499100, 832500000,
    832500900, 832501800, 832502700, 832503600, 832504500, 832505400,
    832506300, 832507200, 832508100, 832509000, 832509900, 832510800,
    832511700, 832512600, 832513500, 832514400, 832515300, 832516200,
    832517100, 832518000, 832518900, 832519800, 832520700, 832521600,
    832522500, 832523400, 832524300, 832525200, 832526100, 832527000,
    832527900, 832528800, 832529700, 832530600, 832531500, 832532400,
    832533300, 832534200, 832535100, 832536000, 832536900, 832537800,
    832538700, 832539600, 832540500, 832541400, 832542300, 832543200,
    832544100, 832545000, 832545900, 832546800, 832547700, 832548600,
    832549500, 832550400, 832551300, 832552200, 832553100, 832554000,
    832554900, 832555800, 832556700, 832557600, 832558500, 832559400,
    832560300, 832561200, 832562100, 832563000, 832563900, 832564800,
    832565700, 832566600, 832567500, 832568400, 832569300, 832570200,
    832571100, 832572000, 832572900, 832573800, 832574700, 832575600,
    832576500, 832577400, 832578300, 832579200, 832580100, 832581000,
    832581900, 832582800, 832583700, 832584600, 832585500, 832586400,
    832587300, 832588200, 832589100, 832590000, 832590900, 832591800,
    832592700, 832593600, 832594500, 832595400, 832596300, 832597200,
    832598100, 832599000, 832599900, 832600800, 832601700, 832602600,
    832603500, 832604400, 832605300, 832606200, 832607100, 832608000,
    832608900, 832609800, 832610700, 832611600, 832612500, 832613400,
    832614300, 832615200, 832616100, 832617000, 832617900, 832618800,
    832619700, 832620600, 832621500, 832622400, 832623300, 832624200,
    832625100, 832626000, 832626900, 832627800, 832628700, 832629600,
    832630500, 832631400, 832632300, 832633200, 832634100, 832635000,
    832635900, 832636800, 832637700, 832638600, 832639500, 832640400,
    832641300, 832642200, 832643100, 832644000, 832644900, 832645800,
    832646700, 832647600, 832648500, 832649400, 832650300, 832651200,
    832652100, 832653000, 832653900, 832654800, 832655700, 832656600,
    832657500, 832658400, 832659300, 832660200, 832661100, 832662000,
    832662900, 832663800, 832664700, 832665600, 832666500, 832667400,
    832668300, 832669200, 832670100, 832671000, 832671900, 832672800,
    832673700, 832674600, 832675500, 832676400, 832677300, 832678200,
    832679100, 832680000, 832680900, 832681800, 832682700, 832683600,
    832684500, 832685400, 832686300, 832687200, 832688100, 832689000,
    832689900, 832690800, 832691700, 832692600, 832693500, 832694400,
    832695300, 832696200, 832697100, 832698000, 832698900, 832699800,
    832700700, 832701600, 832702500, 832703400, 832704300, 832705200,
    832706100, 832707000, 832707900, 832708800, 832709700, 832710600,
    832711500, 832712400, 832713300, 832714200, 832715100, 832716000,
    832716900, 832717800, 832718700, 832719600, 832720500, 832721400,
    832722300, 832723200, 832724100, 832725000, 832725900, 832726800,
    832727700, 832728600, 832729500, 832730400, 832731300, 832732200,
    832733100, 832734000, 832734900, 832735800, 832736700, 832737600,
    832738500, 832739400, 832740300, 832741200, 832742100, 832743000,
    832743900, 832744800, 832745700, 832746600, 832747500, 832748400,
    832749300, 832750200, 832751100, 832752000, 832752900, 832753800,
    832754700, 832755600, 832756500, 832757400, 832758300, 832759200,
    832760100, 832761000, 832761900, 832762800, 832763700, 832764600,
    832765500, 832766400, 832767300, 832768200, 832769100, 832770000,
    832770900, 832771800, 832772700, 832773600, 832774500, 832775400,
    832776300, 832777200, 832778100, 832779000, 832779900, 832780800,
    832781700, 832782600, 832783500, 832784400, 832785300, 832786200,
    832787100, 832788000, 832788900, 832789800, 832790700, 832791600,
    832792500, 832793400, 832794300, 832795200, 832796100, 832797000,
    832797900, 832798800, 832799700, 832800600, 832801500, 832802400,
    832803300, 832804200, 832805100, 832806000, 832806900, 832807800,
    832808700, 832809600, 832810500, 832811400, 832812300, 832813200,
    832814100, 832815000, 832815900, 832816800, 832817700, 832818600,
    832819500, 832820400, 832821300, 832822200, 832823100, 832824000,
    832824900, 832825800, 832826700, 832827600, 832828500, 832829400,
    832830300, 832831200, 832832100, 832833000, 832833900, 832834800,
    832835700, 832836600, 832837500, 832838400, 832839300, 832840200,
    832841100, 832842000, 832842900, 832843800, 832844700, 832845600,
    832846500, 832847400, 832848300, 832849200, 832850100, 832851000,
    832851900, 832852800, 832853700, 832854600, 832855500, 832856400,
    832857300, 832858200, 832859100, 832860000, 832860900, 832861800,
    832862700, 832863600, 832864500, 832865400, 832866300, 832867200,
    832868100, 832869000, 832869900, 832870800, 832871700, 832872600,
    832873500, 832874400, 832875300, 832876200, 832877100, 832878000,
    832878900, 832879800, 832880700, 832881600, 832882500, 832883400,
    832884300, 832885200, 832886100, 832887000, 832887900, 832888800,
    832889700, 832890600, 832891500, 832892400, 832893300, 832894200,
    832895100, 832896000, 832896900, 832897800, 832898700, 832899600,
    832900500, 832901400, 832902300, 832903200, 832904100, 832905000,
    832905900, 832906800, 832907700, 832908600, 832909500, 832910400,
    832911300, 832912200, 832913100, 832914000, 832914900, 832915800,
    832916700, 832917600, 832918500, 832919400, 832920300, 832921200,
    832922100, 832923000, 832923900, 832924800, 832925700, 832926600,
    832927500, 832928400, 832929300, 832930200, 832931100, 832932000,
    832932900, 832933800, 832934700, 832935600, 832936500, 832937400,
    832938300, 832939200, 832940100, 832941000, 832941900, 832942800,
    832943700, 832944600, 832945500, 832946400, 832947300, 832948200,
    832949100, 832950000, 832950900, 832951800, 832952700, 832953600,
    832954500, 832955400, 832956300, 832957200, 832958100, 832959000,
    832959900, 832960800, 832961700, 832962600, 832963500, 832964400,
    832965300, 832966200, 832967100, 832968000, 832968900, 832969800,
    832970700, 832971600, 832972500, 832973400, 832974300, 832975200,
    832976100, 832977000, 832977900, 832978800, 832979700, 832980600,
    832981500, 832982400, 832983300, 832984200, 832985100, 832986000,
    832986900, 832987800, 832988700, 832989600, 832990500, 832991400,
    832992300, 832993200, 832994100, 832995000, 832995900, 832996800,
    832997700, 832998600, 832999500, 833000400, 833001300, 833002200,
    833003100, 833004000, 833004900, 833005800, 833006700, 833007600,
    833008500, 833009400, 833010300, 833011200, 833012100, 833013000,
    833013900, 833014800, 833015700, 833016600, 833017500, 833018400,
    833019300, 833020200, 833021100, 833022000, 833022900, 833023800,
    833024700, 833025600, 833026500, 833027400, 833028300, 833029200,
    833030100, 833031000, 833031900, 833032800, 833033700, 833034600,
    833035500, 833036400, 833037300, 833038200, 833039100, 833040000,
    833040900, 833041800, 833042700, 833043600, 833044500, 833045400,
    833046300, 833047200, 833048100, 833049000, 833049900, 833050800,
    833051700, 833052600, 833053500, 833054400, 833055300, 833056200,
    833057100, 833058000, 833058900, 833059800, 833060700, 833061600,
    833062500, 833063400, 833064300, 833065200, 833066100, 833067000,
    833067900, 833068800, 833069700, 833070600, 833071500, 833072400,
    833073300, 833074200, 833075100, 833076000, 833076900, 833077800,
    833078700, 833079600, 833080500, 833081400, 833082300, 833083200,
    833084100, 833085000, 833085900, 833086800, 833087700, 833088600,
    833089500, 833090400, 833091300, 833092200, 833093100, 833094000,
    833094900, 833095800, 833096700, 833097600, 833098500, 833099400,
    833100300, 833101200, 833102100, 833103000, 833103900, 833104800,
    833105700, 833106600, 833107500, 833108400, 833109300, 833110200,
    833111100, 833112000, 833112900, 833113800, 833114700, 833115600,
    833116500, 833117400, 833118300, 833119200, 833120100, 833121000,
    833121900, 833122800, 833123700, 833124600, 833125500, 833126400,
    833127300, 833128200, 833129100, 833130000, 833130900, 833131800,
    833132700, 833133600, 833134500, 833135400, 833136300, 833137200,
    833138100, 833139000, 833139900, 833140800, 833141700, 833142600,
    833143500, 833144400, 833145300, 833146200, 833147100, 833148000,
    833148900, 833149800, 833150700, 833151600, 833152500, 833153400,
    833154300, 833155200, 833156100, 833157000, 833157900, 833158800,
    833159700, 833160600, 833161500, 833162400, 833163300, 833164200,
    833165100, 833166000, 833166900, 833167800, 833168700, 833169600,
    833170500, 833171400, 833172300, 833173200, 833174100, 833175000,
    833175900, 833176800, 833177700, 833178600, 833179500, 833180400,
    833181300, 833182200, 833183100, 833184000, 833184900, 833185800,
    833186700, 833187600, 833188500, 833189400, 833190300, 833191200,
    833192100, 833193000, 833193900, 833194800, 833195700, 833196600,
    833197500, 833198400, 833199300, 833200200, 833201100, 833202000,
    833202900, 833203800, 833204700, 833205600, 833206500, 833207400,
    833208300, 833209200, 833210100, 833211000, 833211900, 833212800,
    833213700, 833214600, 833215500, 833216400, 833217300, 833218200,
    833219100, 833220000, 833220900, 833221800, 833222700, 833223600,
    833224500, 833225400, 833226300, 833227200, 833228100, 833229000,
    833229900, 833230800, 833231700, 833232600, 833233500, 833234400,
    833235300, 833236200, 833237100, 833238000, 833238900, 833239800,
    833240700, 833241600, 833242500, 833243400, 833244300, 833245200,
    833246100, 833247000, 833247900, 833248800, 833249700, 833250600,
    833251500, 833252400, 833253300, 833254200, 833255100, 833256000,
    833256900, 833257800, 833258700, 833259600, 833260500, 833261400,
    833262300, 833263200, 833264100, 833265000, 833265900, 833266800,
    833267700, 833268600, 833269500, 833270400, 833271300, 833272200,
    833273100, 833274000, 833274900, 833275800, 833276700, 833277600,
    833278500, 833279400, 833280300, 833281200, 833282100, 833283000,
    833283900, 833284800, 833285700, 833286600, 833287500, 833288400,
    833289300, 833290200, 833291100, 833292000, 833292900, 833293800,
    833294700, 833295600, 833296500, 833297400, 833298300, 833299200,
    833300100, 833301000, 833301900, 833302800, 833303700, 833304600,
    833305500, 833306400, 833307300, 833308200, 833309100, 833310000,
    833310900, 833311800, 833312700, 833313600, 833314500, 833315400,
    833316300, 833317200, 833318100, 833319000, 833319900, 833320800,
    833321700, 833322600, 833323500, 833324400, 833325300, 833326200,
    833327100, 833328000, 833328900, 833329800, 833330700, 833331600,
    833332500, 833333400, 833334300, 833335200, 833336100, 833337000,
    833337900, 833338800, 833339700, 833340600, 833341500, 833342400,
    833343300, 833344200, 833345100, 833346000, 833346900, 833347800,
    833348700, 833349600, 833350500, 833351400, 833352300, 833353200,
    833354100, 833355000, 833355900, 833356800, 833357700, 833358600,
    833359500, 833360400, 833361300, 833362200, 833363100, 833364000,
    833364900, 833365800, 833366700, 833367600, 833368500, 833369400,
    833370300, 833371200, 833372100, 833373000, 833373900, 833374800,
    833375700, 833376600, 833377500, 833378400, 833379300, 833380200,
    833381100, 833382000, 833382900, 833383800, 833384700, 833385600,
    833386500, 833387400, 833388300, 833389200, 833390100, 833391000,
    833391900, 833392800, 833393700, 833394600, 833395500, 833396400,
    833397300, 833398200, 833399100, 833400000, 833400900, 833401800,
    833402700, 833403600, 833404500, 833405400, 833406300, 833407200,
    833408100, 833409000, 833409900, 833410800, 833411700, 833412600,
    833413500, 833414400, 833415300, 833416200, 833417100, 833418000,
    833418900, 833419800, 833420700, 833421600, 833422500, 833423400,
    833424300, 833425200, 833426100, 833427000, 833427900, 833428800,
    833429700, 833430600, 833431500, 833432400, 833433300, 833434200,
    833435100, 833436000, 833436900, 833437800, 833438700, 833439600,
    833440500, 833441400, 833442300, 833443200, 833444100, 833445000,
    833445900, 833446800, 833447700, 833448600, 833449500, 833450400,
    833451300, 833452200, 833453100, 833454000, 833454900, 833455800,
    833456700, 833457600, 833458500, 833459400, 833460300, 833461200,
    833462100, 833463000, 833463900, 833464800, 833465700, 833466600,
    833467500, 833468400, 833469300, 833470200, 833471100, 833472000,
    833472900, 833473800, 833474700, 833475600, 833476500, 833477400,
    833478300, 833479200, 833480100, 833481000, 833481900, 833482800,
    833483700, 833484600, 833485500, 833486400, 833487300, 833488200,
    833489100, 833490000, 833490900, 833491800, 833492700, 833493600,
    833494500, 833495400, 833496300, 833497200, 833498100, 833499000,
    833499900, 833500800, 833501700, 833502600, 833503500, 833504400,
    833505300, 833506200, 833507100, 833508000, 833508900, 833509800,
    833510700, 833511600, 833512500, 833513400, 833514300, 833515200,
    833516100, 833517000, 833517900, 833518800, 833519700, 833520600,
    833521500, 833522400, 833523300, 833524200, 833525100, 833526000,
    833526900, 833527800, 833528700, 833529600, 833530500, 833531400,
    833532300, 833533200, 833534100, 833535000, 833535900, 833536800,
    833537700, 833538600, 833539500, 833540400, 833541300, 833542200,
    833543100, 833544000, 833544900, 833545800, 833546700, 833547600,
    833548500, 833549400, 833550300, 833551200, 833552100, 833553000,
    833553900, 833554800, 833555700, 833556600, 833557500, 833558400,
    833559300, 833560200, 833561100, 833562000, 833562900, 833563800,
    833564700, 833565600, 833566500, 833567400, 833568300, 833569200,
    833570100, 833571000, 833571900, 833572800, 833573700, 833574600,
    833575500, 833576400, 833577300, 833578200, 833579100, 833580000,
    833580900, 833581800, 833582700, 833583600, 833584500, 833585400,
    833586300, 833587200, 833588100, 833589000, 833589900, 833590800,
    833591700, 833592600, 833593500, 833594400, 833595300, 833596200,
    833597100, 833598000, 833598900, 833599800, 833600700, 833601600,
    833602500, 833603400, 833604300, 833605200, 833606100, 833607000,
    833607900, 833608800, 833609700, 833610600, 833611500, 833612400,
    833613300, 833614200, 833615100, 833616000, 833616900, 833617800,
    833618700, 833619600, 833620500, 833621400, 833622300, 833623200,
    833624100, 833625000, 833625900, 833626800, 833627700, 833628600,
    833629500, 833630400, 833631300, 833632200, 833633100, 833634000,
    833634900, 833635800, 833636700, 833637600, 833638500, 833639400,
    833640300, 833641200, 833642100, 833643000, 833643900, 833644800,
    833645700, 833646600, 833647500, 833648400, 833649300, 833650200,
    833651100, 833652000, 833652900, 833653800, 833654700, 833655600,
    833656500, 833657400, 833658300, 833659200, 833660100, 833661000,
    833661900, 833662800, 833663700, 833664600, 833665500, 833666400,
    833667300, 833668200, 833669100, 833670000, 833670900, 833671800,
    833672700, 833673600, 833674500, 833675400, 833676300, 833677200,
    833678100, 833679000, 833679900, 833680800, 833681700, 833682600,
    833683500, 833684400, 833685300, 833686200, 833687100, 833688000,
    833688900, 833689800, 833690700, 833691600, 833692500, 833693400,
    833694300, 833695200, 833696100, 833697000, 833697900, 833698800,
    833699700, 833700600, 833701500, 833702400, 833703300, 833704200,
    833705100, 833706000, 833706900, 833707800, 833708700, 833709600,
    833710500, 833711400, 833712300, 833713200, 833714100, 833715000,
    833715900, 833716800, 833717700, 833718600, 833719500, 833720400,
    833721300, 833722200, 833723100, 833724000, 833724900, 833725800,
    833726700, 833727600, 833728500, 833729400, 833730300, 833731200,
    833732100, 833733000, 833733900, 833734800, 833735700, 833736600,
    833737500, 833738400, 833739300, 833740200, 833741100, 833742000,
    833742900, 833743800, 833744700, 833745600, 833746500, 833747400,
    833748300, 833749200, 833750100, 833751000, 833751900, 833752800,
    833753700, 833754600, 833755500, 833756400, 833757300, 833758200,
    833759100, 833760000, 833760900, 833761800, 833762700, 833763600,
    833764500, 833765400, 833766300, 833767200, 833768100, 833769000,
    833769900, 833770800, 833771700, 833772600, 833773500, 833774400,
    833775300, 833776200, 833777100, 833778000, 833778900, 833779800,
    833780700, 833781600, 833782500, 833783400, 833784300, 833785200,
    833786100, 833787000, 833787900, 833788800, 833789700, 833790600,
    833791500, 833792400, 833793300, 833794200, 833795100, 833796000,
    833796900, 833797800, 833798700, 833799600, 833800500, 833801400,
    833802300, 833803200, 833804100, 833805000, 833805900, 833806800,
    833807700, 833808600, 833809500, 833810400, 833811300, 833812200,
    833813100, 833814000, 833814900, 833815800, 833816700, 833817600,
    833818500, 833819400, 833820300, 833821200, 833822100, 833823000,
    833823900, 833824800, 833825700, 833826600, 833827500, 833828400,
    833829300, 833830200, 833831100, 833832000, 833832900, 833833800,
    833834700, 833835600, 833836500, 833837400, 833838300, 833839200,
    833840100, 833841000, 833841900, 833842800, 833843700, 833844600,
    833845500, 833846400, 833847300, 833848200, 833849100, 833850000,
    833850900, 833851800, 833852700, 833853600, 833854500, 833855400,
    833856300, 833857200, 833858100, 833859000, 833859900, 833860800,
    833861700, 833862600, 833863500, 833864400, 833865300, 833866200,
    833867100, 833868000, 833868900, 833869800, 833870700, 833871600,
    833872500, 833873400, 833874300, 833875200, 833876100, 833877000,
    833877900, 833878800, 833879700, 833880600, 833881500, 833882400,
    833883300, 833884200, 833885100, 833886000, 833886900, 833887800,
    833888700, 833889600, 833890500, 833891400, 833892300, 833893200,
    833894100, 833895000, 833895900, 833896800, 833897700, 833898600,
    833899500, 833900400, 833901300, 833902200, 833903100, 833904000,
    833904900, 833905800, 833906700, 833907600, 833908500, 833909400,
    833910300, 833911200, 833912100, 833913000, 833913900, 833914800,
    833915700, 833916600, 833917500, 833918400, 833919300, 833920200,
    833921100, 833922000, 833922900, 833923800, 833924700, 833925600,
    833926500, 833927400, 833928300, 833929200, 833930100, 833931000,
    833931900, 833932800, 833933700, 833934600, 833935500, 833936400,
    833937300, 833938200, 833939100, 833940000, 833940900, 833941800,
    833942700, 833943600, 833944500, 833945400, 833946300, 833947200,
    833948100, 833949000, 833949900, 833950800, 833951700, 833952600,
    833953500, 833954400, 833955300, 833956200, 833957100, 833958000,
    833958900, 833959800, 833960700, 833961600, 833962500, 833963400,
    833964300, 833965200, 833966100, 833967000, 833967900, 833968800,
    833969700, 833970600, 833971500, 833972400, 833973300, 833974200,
    833975100, 833976000, 833976900, 833977800, 833978700, 833979600,
    833980500, 833981400, 833982300, 833983200, 833984100, 833985000,
    833985900, 833986800, 833987700, 833988600, 833989500, 833990400,
    833991300, 833992200, 833993100, 833994000, 833994900, 833995800,
    833996700, 833997600, 833998500, 833999400, 834000300, 834001200,
    834002100, 834003000, 834003900, 834004800, 834005700, 834006600,
    834007500, 834008400, 834009300, 834010200, 834011100, 834012000,
    834012900, 834013800, 834014700, 834015600, 834016500, 834017400,
    834018300, 834019200, 834020100, 834021000, 834021900, 834022800,
    834023700, 834024600, 834025500, 834026400, 834027300, 834028200,
    834029100, 834030000, 834030900, 834031800, 834032700, 834033600,
    834034500, 834035400, 834036300, 834037200, 834038100, 834039000,
    834039900, 834040800, 834041700, 834042600, 834043500, 834044400,
    834045300, 834046200, 834047100, 834048000, 834048900, 834049800,
    834050700, 834051600, 834052500, 834053400, 834054300, 834055200,
    834056100, 834057000, 834057900, 834058800, 834059700, 834060600,
    834061500, 834062400, 834063300, 834064200, 834065100, 834066000,
    834066900, 834067800, 834068700, 834069600, 834070500, 834071400,
    834072300, 834073200, 834074100, 834075000, 834075900, 834076800,
    834077700, 834078600, 834079500, 834080400, 834081300, 834082200,
    834083100, 834084000, 834084900, 834085800, 834086700, 834087600,
    834088500, 834089400, 834090300, 834091200, 834092100, 834093000,
    834093900, 834094800, 834095700, 834096600, 834097500, 834098400,
    834099300, 834100200, 834101100, 834102000, 834102900, 834103800,
    834104700, 834105600, 834106500, 834107400, 834108300, 834109200,
    834110100, 834111000, 834111900, 834112800, 834113700, 834114600,
    834115500, 834116400, 834117300, 834118200, 834119100, 834120000,
    834120900, 834121800, 834122700, 834123600, 834124500, 834125400,
    834126300, 834127200, 834128100, 834129000, 834129900, 834130800,
    834131700, 834132600, 834133500, 834134400, 834135300, 834136200,
    834137100, 834138000, 834138900, 834139800, 834140700, 834141600,
    834142500, 834143400, 834144300, 834145200, 834146100, 834147000,
    834147900, 834148800, 834149700, 834150600, 834151500, 834152400,
    834153300, 834154200, 834155100, 834156000, 834156900, 834157800,
    834158700, 834159600, 834160500, 834161400, 834162300, 834163200,
    834164100, 834165000, 834165900, 834166800, 834167700, 834168600,
    834169500, 834170400, 834171300, 834172200, 834173100, 834174000,
    834174900, 834175800, 834176700, 834177600, 834178500, 834179400,
    834180300, 834181200, 834182100, 834183000, 834183900, 834184800,
    834185700, 834186600, 834187500, 834188400, 834189300, 834190200,
    834191100, 834192000, 834192900, 834193800, 834194700, 834195600,
    834196500, 834197400, 834198300, 834199200, 834200100, 834201000,
    834201900, 834202800, 834203700, 834204600, 834205500, 834206400,
    834207300, 834208200, 834209100, 834210000, 834210900, 834211800,
    834212700, 834213600, 834214500, 834215400, 834216300, 834217200,
    834218100, 834219000, 834219900, 834220800, 834221700, 834222600,
    834223500, 834224400, 834225300, 834226200, 834227100, 834228000,
    834228900, 834229800, 834230700, 834231600, 834232500, 834233400,
    834234300, 834235200, 834236100, 834237000, 834237900, 834238800,
    834239700, 834240600, 834241500, 834242400, 834243300, 834244200,
    834245100, 834246000, 834246900, 834247800, 834248700, 834249600,
    834250500, 834251400, 834252300, 834253200, 834254100, 834255000,
    834255900, 834256800, 834257700, 834258600, 834259500, 834260400,
    834263100, 834264000, 834264900, 834265800, 834266700, 834267600,
    834268500, 834269400, 834270300, 834271200, 834272100, 834273000,
    834273900, 834274800, 834275700, 834276600, 834277500, 834278400,
    834279300, 834280200, 834281100, 834282000, 834282900, 834283800,
    834284700, 834285600, 834286500, 834287400, 834288300, 834289200,
    834290100, 834291000, 834291900, 834292800, 834293700, 834294600,
    834295500, 834296400, 834297300, 834298200, 834299100, 834300000,
    834300900, 834301800, 834302700, 834303600, 834304500, 834305400,
    834306300, 834307200, 834308100, 834309000, 834309900, 834310800,
    834311700, 834312600, 834313500, 834314400, 834315300, 834316200,
    834317100, 834318000, 834318900, 834319800, 834320700, 834321600,
    834322500, 834323400, 834324300, 834325200, 834326100, 834327000,
    834327900, 834328800, 834329700, 834330600, 834331500, 834332400,
    834333300, 834334200, 834335100, 834336000, 834336900, 834337800,
    834338700, 834339600, 834340500, 834341400, 834342300, 834343200,
    834344100, 834345000, 834345900, 834346800, 834347700, 834348600,
    834349500, 834350400, 834351300, 834352200, 834353100, 834354000,
    834354900, 834355800, 834356700, 834357600, 834358500, 834359400,
    834360300, 834361200, 834362100, 834363000, 834363900, 834364800,
    834365700, 834366600, 834367500, 834368400, 834369300, 834370200,
    834371100, 834372000, 834372900, 834373800, 834374700, 834375600,
    834376500, 834377400, 834378300, 834379200, 834380100, 834381000,
    834381900, 834382800, 834383700, 834384600, 834385500, 834386400,
    834387300, 834388200, 834389100, 834390000, 834390900, 834391800,
    834392700, 834393600, 834394500, 834395400, 834396300, 834397200,
    834398100, 834399000, 834399900, 834400800, 834401700, 834402600,
    834403500, 834404400, 834405300, 834406200, 834407100, 834408000,
    834408900, 834409800, 834410700, 834411600, 834412500, 834413400,
    834414300, 834415200, 834416100, 834417000, 834417900, 834418800,
    834419700, 834420600, 834421500, 834422400, 834423300, 834424200,
    834425100, 834426000, 834426900, 834427800, 834428700, 834429600,
    834430500, 834431400, 834432300, 834433200, 834434100, 834435000,
    834435900, 834436800, 834437700, 834438600, 834439500, 834440400,
    834441300, 834442200, 834443100, 834444000, 834444900, 834445800,
    834446700, 834447600, 834448500, 834449400, 834450300, 834451200,
    834452100, 834453000, 834453900, 834454800, 834455700, 834456600,
    834457500, 834458400, 834459300, 834460200, 834461100, 834462000,
    834462900, 834463800, 834464700, 834465600, 834466500, 834467400,
    834468300, 834469200, 834470100, 834471000, 834471900, 834472800,
    834473700, 834474600, 834475500, 834476400, 834477300, 834478200,
    834479100, 834480000, 834480900, 834481800, 834482700, 834483600,
    834484500, 834485400, 834486300, 834487200, 834488100, 834489000,
    834489900, 834490800, 834491700, 834492600, 834493500, 834494400,
    834495300, 834496200, 834497100, 834498000, 834498900, 834499800,
    834500700, 834501600, 834502500, 834503400, 834504300, 834505200,
    834506100, 834507000, 834507900, 834508800, 834509700, 834510600,
    834511500, 834512400, 834513300, 834514200, 834515100, 834516000,
    834516900, 834517800, 834518700, 834519600, 834520500, 834521400,
    834522300, 834523200, 834524100, 834525000, 834525900, 834526800,
    834527700, 834528600, 834529500, 834530400, 834531300, 834532200,
    834533100, 834534000, 834534900, 834535800, 834536700, 834537600,
    834538500, 834539400, 834540300, 834541200, 834542100, 834543000,
    834543900, 834544800, 834545700, 834546600, 834547500, 834548400,
    834549300, 834550200, 834551100, 834552000, 834552900, 834553800,
    834554700, 834555600, 834556500, 834557400, 834558300, 834559200,
    834560100, 834561000, 834561900, 834562800, 834563700, 834564600,
    834565500, 834566400, 834567300, 834568200, 834569100, 834570000,
    834570900, 834571800, 834572700, 834573600, 834574500, 834575400,
    834576300, 834577200, 834578100, 834579000, 834579900, 834580800,
    834581700, 834582600, 834583500, 834584400, 834585300, 834586200,
    834587100, 834588000, 834588900, 834589800, 834590700, 834591600,
    834592500, 834593400, 834594300, 834595200, 834596100, 834597000,
    834597900, 834598800, 834599700, 834600600, 834601500, 834602400,
    834603300, 834604200, 834605100, 834606000, 834606900, 834607800,
    834608700, 834609600, 834610500, 834611400, 834612300, 834613200,
    834614100, 834615000, 834615900, 834616800, 834617700, 834618600,
    834619500, 834620400, 834621300, 834622200, 834623100, 834624000,
    834624900, 834625800, 834626700, 834627600, 834628500, 834629400,
    834630300, 834631200, 834632100, 834633000, 834633900, 834634800,
    834635700, 834636600, 834637500, 834638400, 834639300, 834640200,
    834641100, 834642000, 834642900, 834643800, 834644700, 834645600,
    834646500, 834647400, 834648300, 834649200, 834650100, 834651000,
    834651900, 834652800, 834653700, 834654600, 834655500, 834656400,
    834657300, 834658200, 834659100, 834660000, 834660900, 834661800,
    834662700, 834663600, 834664500, 834665400, 834666300, 834667200,
    834668100, 834669000, 834669900, 834670800, 834671700, 834672600,
    834673500, 834674400, 834675300, 834676200, 834677100, 834678000,
    834678900, 834679800, 834680700, 834681600, 834682500, 834683400,
    834684300, 834685200, 834686100, 834687000, 834687900, 834688800,
    834689700, 834690600, 834691500, 834692400, 834693300, 834694200,
    834695100, 834696000, 834696900, 834697800, 834698700, 834699600,
    834700500, 834701400, 834702300, 834703200, 834704100, 834705000,
    834705900, 834706800, 834707700, 834708600, 834709500, 834710400,
    834711300, 834712200, 834713100, 834714000, 834714900, 834715800,
    834716700, 834717600, 834718500, 834719400, 834720300, 834721200,
    834722100, 834723000, 834723900, 834724800, 834725700, 834726600,
    834727500, 834728400, 834729300, 834730200, 834731100, 834732000,
    834732900, 834733800, 834734700, 834735600, 834736500, 834737400,
    834738300, 834739200, 834740100, 834741000, 834741900, 834742800,
    834743700, 834744600, 834745500, 834746400, 834747300, 834748200,
    834749100, 834750000, 834750900, 834751800, 834752700, 834753600,
    834754500, 834755400, 834756300, 834757200, 834758100, 834759000,
    834759900, 834760800, 834761700, 834762600, 834763500, 834764400,
    834765300, 834766200, 834767100, 834768000, 834768900, 834769800,
    834770700, 834771600, 834772500, 834773400, 834774300, 834775200,
    834776100, 834777000, 834777900, 834778800, 834779700, 834780600,
    834781500, 834782400, 834783300, 834784200, 834785100, 834786000,
    834786900, 834787800, 834788700, 834789600, 834790500, 834791400,
    834792300, 834793200, 834794100, 834795000, 834795900, 834796800,
    834797700, 834798600, 834799500, 834800400, 834801300, 834802200,
    834803100, 834804000, 834804900, 834805800, 834806700, 834807600,
    834808500, 834809400, 834810300, 834811200, 834812100, 834813000,
    834813900, 834814800, 834815700, 834816600, 834817500, 834818400,
    834819300, 834820200, 834821100, 834822000, 834822900, 834823800,
    834824700, 834825600, 834826500, 834827400, 834828300, 834829200,
    834830100, 834831000, 834831900, 834832800, 834833700, 834834600,
    834835500, 834836400, 834837300, 834838200, 834839100, 834840000,
    834840900, 834841800, 834842700, 834843600, 834844500, 834845400,
    834846300, 834847200, 834848100, 834849000, 834849900, 834850800,
    834851700, 834852600, 834853500, 834854400, 834855300, 834856200,
    834857100, 834858000, 834858900, 834859800, 834860700, 834861600,
    834862500, 834863400, 834864300, 834865200, 834866100, 834867000,
    834867900, 834868800, 834869700, 834870600, 834871500, 834872400,
    834873300, 834874200, 834875100, 834876000, 834876900, 834877800,
    834878700, 834879600, 834880500, 834881400, 834882300, 834883200,
    834884100, 834885000, 834885900, 834886800, 834887700, 834888600,
    834889500, 834890400, 834891300, 834892200, 834893100, 834894000,
    834894900, 834895800, 834896700, 834897600, 834898500, 834899400,
    834900300, 834901200, 834902100, 834903000, 834903900, 834904800,
    834905700, 834906600, 834907500, 834908400, 834909300, 834910200,
    834911100, 834912000, 834912900, 834913800, 834914700, 834915600,
    834916500, 834917400, 834918300, 834919200, 834920100, 834921000,
    834921900, 834922800, 834923700, 834924600, 834925500, 834926400,
    834927300, 834928200, 834929100, 834930000, 834930900, 834931800,
    834932700, 834933600, 834934500, 834935400, 834936300, 834937200,
    834938100, 834939000, 834939900, 834940800, 834941700, 834942600,
    834943500, 834944400, 834945300, 834946200, 834947100, 834948000,
    834948900, 834949800, 834950700, 834951600, 834952500, 834953400,
    834954300, 834955200, 834956100, 834957000, 834957900, 834958800,
    834959700, 834960600, 834961500, 834962400, 834963300, 834964200,
    834965100, 834966000, 834966900, 834967800, 834968700, 834969600,
    834970500, 834971400, 834972300, 834973200, 834974100, 834975000,
    834975900, 834976800, 834977700, 834978600, 834979500, 834980400,
    834981300, 834982200, 834983100, 834984000, 834984900, 834985800,
    834986700, 834987600, 834988500, 834989400, 834990300, 834991200,
    834992100, 834993000, 834993900, 834994800, 834995700, 834996600,
    834997500, 834998400, 834999300, 835000200, 835001100, 835002000,
    835002900, 835003800, 835004700, 835005600, 835006500, 835007400,
    835008300, 835009200, 835010100, 835011000, 835011900, 835012800,
    835013700, 835014600, 835015500, 835016400, 835017300, 835018200,
    835019100, 835020000, 835020900, 835021800, 835022700, 835023600,
    835024500, 835025400, 835026300, 835027200, 835028100, 835029000,
    835029900, 835030800, 835031700, 835032600, 835033500, 835034400,
    835035300, 835036200, 835037100, 835038000, 835038900, 835039800,
    835040700, 835041600, 835042500, 835043400, 835044300, 835045200,
    835046100, 835047000, 835047900, 835048800, 835049700, 835050600,
    835051500, 835052400, 835053300, 835054200, 835055100, 835056000,
    835056900, 835057800, 835058700, 835059600, 835060500, 835061400,
    835062300, 835063200, 835064100, 835065000, 835065900, 835066800,
    835067700, 835068600, 835069500, 835070400, 835071300, 835072200,
    835073100, 835074000, 835074900, 835075800, 835076700, 835077600,
    835078500, 835079400, 835080300, 835081200, 835082100, 835083000,
    835083900, 835084800, 835085700, 835086600, 835087500, 835088400,
    835089300, 835090200, 835091100, 835092000, 835092900, 835093800,
    835094700, 835095600, 835096500, 835097400, 835098300, 835099200,
    835100100, 835101000, 835101900, 835102800, 835103700, 835104600,
    835105500, 835106400, 835107300, 835108200, 835109100, 835110000,
    835110900, 835111800, 835112700, 835113600, 835114500, 835115400,
    835116300, 835117200, 835118100, 835119000, 835119900, 835120800,
    835121700, 835122600, 835123500, 835124400, 835125300, 835126200,
    835127100, 835128000, 835128900, 835129800, 835130700, 835131600,
    835132500, 835133400, 835134300, 835135200, 835136100, 835137000,
    835137900, 835138800, 835139700, 835140600, 835141500, 835142400,
    835143300, 835144200, 835145100, 835146000, 835146900, 835147800,
    835148700, 835149600, 835150500, 835151400, 835152300, 835153200,
    835154100, 835155000, 835155900, 835156800, 835157700, 835158600,
    835159500, 835160400, 835161300, 835162200, 835163100, 835164000,
    835164900, 835165800, 835166700, 835167600, 835168500, 835169400,
    835170300, 835171200, 835172100, 835173000, 835173900, 835174800,
    835175700, 835176600, 835177500, 835178400, 835179300, 835180200,
    835181100, 835182000, 835182900, 835183800, 835184700, 835185600,
    835186500, 835187400, 835188300, 835189200, 835190100, 835191000,
    835191900, 835192800, 835193700, 835194600, 835195500, 835196400,
    835197300, 835198200, 835199100, 835200000, 835200900, 835201800,
    835202700, 835203600, 835204500, 835205400, 835206300, 835207200,
    835208100, 835209000, 835209900, 835210800, 835211700, 835212600,
    835213500, 835214400, 835215300, 835216200, 835217100, 835218000,
    835218900, 835219800, 835220700, 835221600, 835222500, 835223400,
    835224300, 835225200, 835226100, 835227000, 835227900, 835228800,
    835229700, 835230600, 835231500, 835232400, 835233300, 835234200,
    835235100, 835236000, 835236900, 835237800, 835238700, 835239600,
    835240500, 835241400, 835242300, 835243200, 835244100, 835245000,
    835245900, 835246800, 835247700, 835248600, 835249500, 835250400,
    835251300, 835252200, 835253100, 835254000, 835254900, 835255800,
    835256700, 835257600, 835258500, 835259400, 835260300, 835261200,
    835262100, 835263000, 835263900, 835264800, 835265700, 835266600,
    835267500, 835268400, 835269300, 835270200, 835271100, 835272000,
    835272900, 835273800, 835274700, 835275600, 835276500, 835277400,
    835278300, 835279200, 835280100, 835281000, 835281900, 835282800,
    835283700, 835284600, 835285500, 835286400, 835287300, 835288200,
    835289100, 835290000, 835290900, 835291800, 835292700, 835293600,
    835294500, 835295400, 835296300, 835297200, 835298100, 835299000,
    835299900, 835300800, 835301700, 835302600, 835303500, 835304400,
    835305300, 835306200, 835307100, 835308000, 835308900, 835309800,
    835310700, 835311600, 835312500, 835313400, 835314300, 835315200,
    835316100, 835317000, 835317900, 835318800, 835319700, 835320600,
    835321500, 835322400, 835323300, 835324200, 835325100, 835326000,
    835326900, 835327800, 835328700, 835329600, 835330500, 835331400,
    835332300, 835333200, 835334100, 835335000, 835335900, 835336800,
    835337700, 835338600, 835339500, 835340400, 835341300, 835342200,
    835343100, 835344000, 835344900, 835345800, 835346700, 835347600,
    835348500, 835349400, 835350300, 835351200, 835352100, 835353000,
    835353900, 835354800, 835355700, 835356600, 835357500, 835358400,
    835359300, 835360200, 835361100, 835362000, 835362900, 835363800,
    835364700, 835365600, 835366500, 835367400, 835368300, 835369200,
    835370100, 835371000, 835371900, 835372800, 835373700, 835374600,
    835375500, 835376400, 835377300, 835378200, 835379100, 835380000,
    835380900, 835381800, 835382700, 835383600, 835384500, 835385400,
    835386300, 835387200, 835388100, 835389000, 835389900, 835390800,
    835391700, 835392600, 835393500, 835394400, 835395300, 835396200,
    835397100, 835398000, 835398900, 835399800, 835400700, 835401600,
    835402500, 835403400, 835404300, 835405200, 835406100, 835407000,
    835407900, 835408800, 835409700, 835410600, 835411500, 835412400,
    835413300, 835414200, 835415100, 835416000, 835416900, 835417800,
    835418700, 835419600, 835420500, 835421400, 835422300, 835423200,
    835424100, 835425000, 835425900, 835426800, 835427700, 835428600,
    835429500, 835430400, 835431300, 835432200, 835433100, 835434000,
    835434900, 835435800, 835436700, 835437600, 835438500, 835439400,
    835440300, 835441200, 835442100, 835443000, 835443900, 835444800,
    835445700, 835446600, 835447500, 835448400, 835449300, 835450200,
    835451100, 835452000, 835452900, 835453800, 835454700, 835455600,
    835456500, 835457400, 835458300, 835459200, 835460100, 835461000,
    835461900, 835462800, 835463700, 835464600, 835465500, 835466400,
    835467300, 835468200, 835469100, 835470000, 835470900, 835471800,
    835472700, 835473600, 835474500, 835475400, 835476300, 835477200,
    835478100, 835479000, 835479900, 835480800, 835481700, 835482600,
    835483500, 835484400, 835485300, 835486200, 835487100, 835488000,
    835488900, 835489800, 835490700, 835491600, 835492500, 835493400,
    835494300, 835495200, 835496100, 835497000, 835497900, 835498800,
    835499700, 835500600, 835501500, 835502400, 835503300, 835504200,
    835505100, 835506000, 835506900, 835507800, 835508700, 835509600,
    835510500, 835511400, 835512300, 835513200, 835514100, 835515000,
    835515900, 835516800, 835517700, 835518600, 835519500, 835520400,
    835521300, 835522200, 835523100, 835524000, 835524900, 835525800,
    835526700, 835527600, 835528500, 835529400, 835530300, 835531200,
    835532100, 835533000, 835533900, 835534800, 835535700, 835536600,
    835537500, 835538400, 835539300, 835540200, 835541100, 835542000,
    835542900, 835543800, 835544700, 835545600, 835546500, 835547400,
    835548300, 835549200, 835550100, 835551000, 835551900, 835552800,
    835553700, 835554600, 835555500, 835556400, 835557300, 835558200,
    835559100, 835560000, 835560900, 835561800, 835562700, 835563600,
    835564500, 835565400, 835566300, 835567200, 835568100, 835569000,
    835569900, 835570800, 835571700, 835572600, 835573500, 835574400,
    835575300, 835576200, 835577100, 835578000, 835578900, 835579800,
    835580700, 835581600, 835582500, 835583400, 835584300, 835585200,
    835586100, 835587000, 835587900, 835588800, 835589700, 835590600,
    835591500, 835592400, 835593300, 835594200, 835595100, 835596000,
    835596900, 835597800, 835598700, 835599600, 835600500, 835601400,
    835602300, 835603200, 835604100, 835605000, 835605900, 835606800,
    835607700, 835608600, 835609500, 835610400, 835611300, 835612200,
    835613100, 835614000, 835614900, 835615800, 835616700, 835617600,
    835618500, 835619400, 835620300, 835621200, 835622100, 835623000,
    835623900, 835624800, 835625700, 835626600, 835627500, 835628400,
    835629300, 835630200, 835631100, 835632000, 835632900, 835633800,
    835634700, 835635600, 835636500, 835637400, 835638300, 835639200,
    835640100, 835641000, 835641900, 835642800, 835643700, 835644600,
    835645500, 835646400, 835647300, 835648200, 835649100, 835650000,
    835650900, 835651800, 835652700, 835653600, 835654500, 835655400,
    835656300, 835657200, 835658100, 835659000, 835659900, 835660800,
    835661700, 835662600, 835663500, 835664400, 835665300, 835666200,
    835667100, 835668000, 835668900, 835669800, 835670700, 835671600,
    835672500, 835673400, 835674300, 835675200, 835676100, 835677000,
    835677900, 835678800, 835679700, 835680600, 835681500, 835682400,
    835683300, 835684200, 835685100, 835686000, 835686900, 835687800,
    835688700, 835689600, 835690500, 835691400, 835692300, 835693200,
    835694100, 835695000, 835695900, 835696800, 835697700, 835698600,
    835699500, 835700400, 835701300, 835702200, 835703100, 835704000,
    835704900, 835705800, 835706700, 835707600, 835708500, 835709400,
    835710300, 835711200, 835712100, 835713000, 835713900, 835714800,
    835715700, 835716600, 835717500, 835718400, 835719300, 835720200,
    835721100, 835722000, 835722900, 835723800, 835724700, 835725600,
    835726500, 835727400, 835728300, 835729200, 835730100, 835731000,
    835731900, 835732800, 835733700, 835734600, 835735500, 835736400,
    835737300, 835738200, 835739100, 835740000, 835740900, 835741800,
    835742700, 835743600, 835744500, 835745400, 835746300, 835747200,
    835748100, 835749000, 835749900, 835750800, 835751700, 835752600,
    835753500, 835754400, 835755300, 835756200, 835757100, 835758000,
    835758900, 835759800, 835760700, 835761600, 835762500, 835763400,
    835764300, 835765200, 835766100, 835767000, 835767900, 835768800,
    835769700, 835770600, 835771500, 835772400, 835773300, 835774200,
    835775100, 835776000, 835776900, 835777800, 835778700, 835779600,
    835780500, 835781400, 835782300, 835783200, 835784100, 835785000,
    835785900, 835786800, 835787700, 835788600, 835789500, 835790400,
    835791300, 835792200, 835793100, 835794000, 835794900, 835795800,
    835796700, 835797600, 835798500, 835799400, 835800300, 835801200,
    835802100, 835803000, 835803900, 835804800, 835805700, 835806600,
    835807500, 835808400, 835809300, 835810200, 835811100, 835812000,
    835812900, 835813800, 835814700, 835815600, 835816500, 835817400,
    835818300, 835819200, 835820100, 835821000, 835821900, 835822800,
    835823700, 835824600, 835825500, 835826400, 835827300, 835828200,
    835829100, 835830000, 835830900, 835831800, 835832700, 835833600,
    835834500, 835835400, 835836300, 835837200, 835838100, 835839000,
    835839900, 835840800, 835841700, 835842600, 835843500, 835844400,
    835845300, 835846200, 835847100, 835848000, 835848900, 835849800,
    835850700, 835851600, 835852500, 835853400, 835854300, 835855200,
    835856100, 835857000, 835857900, 835858800, 835859700, 835860600,
    835861500, 835862400, 835863300, 835864200, 835865100, 835866000,
    835866900, 835867800, 835868700, 835869600, 835870500, 835871400,
    835872300, 835873200, 835874100, 835875000, 835875900, 835876800,
    835877700, 835878600, 835879500, 835880400, 835881300, 835882200,
    835883100, 835884000, 835884900, 835885800, 835886700, 835887600,
    835888500, 835889400, 835890300, 835891200, 835892100, 835893000,
    835893900, 835894800, 835895700, 835896600, 835897500, 835898400,
    835899300, 835900200, 835901100, 835902000, 835902900, 835903800,
    835904700, 835905600, 835906500, 835907400, 835908300, 835909200,
    835910100, 835911000, 835911900, 835912800, 835913700, 835914600,
    835915500, 835916400, 835917300, 835918200, 835919100, 835920000,
    835920900, 835921800, 835922700, 835923600, 835924500, 835925400,
    835926300, 835927200, 835928100, 835929000, 835929900, 835930800,
    835931700, 835932600, 835933500, 835934400, 835935300, 835936200,
    835937100, 835938000, 835938900, 835939800, 835940700, 835941600,
    835942500, 835943400, 835944300, 835945200, 835946100, 835947000,
    835947900, 835948800, 835949700, 835950600, 835951500, 835952400,
    835953300, 835954200, 835955100, 835956000, 835956900, 835957800,
    835958700, 835959600, 835960500, 835961400, 835962300, 835963200,
    835964100, 835965000, 835965900, 835966800, 835967700, 835968600,
    835969500, 835970400, 835971300, 835972200, 835973100, 835974000,
    835974900, 835975800, 835976700, 835977600, 835978500, 835979400,
    835980300, 835981200, 835982100, 835983000, 835983900, 835984800,
    835985700, 835986600, 835987500, 835988400, 835989300, 835990200,
    835991100, 835992000, 835992900, 835993800, 835994700, 835995600,
    835996500, 835997400, 835998300, 835999200, 836000100, 836001000,
    836001900, 836002800, 836003700, 836004600, 836005500, 836006400,
    836007300, 836008200, 836009100, 836010000, 836010900, 836011800,
    836012700, 836013600, 836014500, 836015400, 836016300, 836017200,
    836018100, 836019000, 836019900, 836020800, 836021700, 836022600,
    836023500, 836024400, 836025300, 836026200, 836027100, 836028000,
    836028900, 836029800, 836030700, 836031600, 836032500, 836033400,
    836034300, 836035200, 836036100, 836037000, 836037900, 836038800,
    836039700, 836040600, 836041500, 836042400, 836043300, 836044200,
    836045100, 836046000, 836046900, 836047800, 836048700, 836049600,
    836050500, 836051400, 836052300, 836053200, 836054100, 836055000,
    836055900, 836056800, 836057700, 836058600, 836059500, 836060400,
    836061300, 836062200, 836063100, 836064000, 836064900, 836065800,
    836066700, 836067600, 836068500, 836069400, 836070300, 836071200,
    836072100, 836073000, 836073900, 836074800, 836075700, 836076600,
    836077500, 836078400, 836079300, 836080200, 836081100, 836082000,
    836082900, 836083800, 836084700, 836085600, 836086500, 836087400,
    836088300, 836089200, 836090100, 836091000, 836091900, 836092800,
    836093700, 836094600, 836095500, 836096400, 836097300, 836098200,
    836099100, 836100000, 836100900, 836101800, 836102700, 836103600,
    836104500, 836105400, 836106300, 836107200, 836108100, 836109000,
    836109900, 836110800, 836111700, 836112600, 836113500, 836114400,
    836115300, 836116200, 836117100, 836118000, 836118900, 836119800,
    836120700, 836121600, 836122500, 836123400, 836124300, 836125200,
    836126100, 836127000, 836127900, 836128800, 836129700, 836130600,
    836131500, 836132400, 836133300, 836134200, 836135100, 836136000,
    836136900, 836137800, 836138700, 836139600, 836140500, 836141400,
    836142300, 836143200, 836144100, 836145000, 836145900, 836146800,
    836147700, 836148600, 836149500, 836150400, 836151300, 836152200,
    836153100, 836154000, 836154900, 836155800, 836156700, 836157600,
    836158500, 836159400, 836160300, 836161200, 836162100, 836163000,
    836163900, 836164800, 836165700, 836166600, 836167500, 836168400,
    836169300, 836170200, 836171100, 836172000, 836172900, 836173800,
    836174700, 836175600, 836176500, 836177400, 836178300, 836179200,
    836180100, 836181000, 836181900, 836182800, 836183700, 836184600,
    836185500, 836186400, 836187300, 836188200, 836189100, 836190000,
    836190900, 836191800, 836192700, 836193600, 836194500, 836195400,
    836196300, 836197200, 836198100, 836199000, 836199900, 836200800,
    836201700, 836202600, 836203500, 836204400, 836205300, 836206200,
    836207100, 836208000, 836208900, 836209800, 836210700, 836211600,
    836212500, 836213400, 836214300, 836215200, 836216100, 836217000,
    836217900, 836218800, 836219700, 836220600, 836221500, 836222400,
    836223300, 836224200, 836225100, 836226000, 836226900, 836227800,
    836228700, 836229600, 836230500, 836231400, 836232300, 836233200,
    836234100, 836235000, 836235900, 836236800, 836239500, 836240400,
    836241300, 836242200, 836243100, 836244000, 836244900, 836245800,
    836246700, 836247600, 836248500, 836249400, 836250300, 836251200,
    836252100, 836253000, 836253900, 836254800, 836255700, 836256600,
    836257500, 836258400, 836259300, 836260200, 836261100, 836262000,
    836262900, 836263800, 836264700, 836265600, 836266500, 836267400,
    836268300, 836269200, 836270100, 836271000, 836271900, 836272800,
    836273700, 836274600, 836275500, 836276400, 836277300, 836278200,
    836279100, 836280000, 836280900, 836281800, 836282700, 836283600,
    836284500, 836285400, 836286300, 836287200, 836288100, 836289000,
    836289900, 836290800, 836291700, 836292600, 836293500, 836294400,
    836295300, 836296200, 836297100, 836298000, 836298900, 836299800,
    836300700, 836301600, 836302500, 836303400, 836304300, 836305200,
    836306100, 836307000, 836307900, 836308800, 836309700, 836310600,
    836311500, 836312400, 836313300, 836314200, 836315100, 836316000,
    836316900, 836317800, 836318700, 836319600, 836320500, 836321400,
    836322300, 836323200, 836324100, 836325000, 836325900, 836326800,
    836327700, 836328600, 836329500, 836330400, 836331300, 836332200,
    836333100, 836334000, 836334900, 836335800, 836336700, 836337600,
    836338500, 836339400, 836340300, 836341200, 836342100, 836343000,
    836343900, 836344800, 836345700, 836346600, 836347500, 836348400,
    836349300, 836350200, 836351100, 836352000, 836352900, 836353800,
    836354700, 836355600, 836356500, 836357400, 836358300, 836359200,
    836360100, 836361000, 836361900, 836362800, 836363700, 836364600,
    836365500, 836366400, 836367300, 836368200, 836369100, 836370000,
    836370900, 836371800, 836372700, 836373600, 836374500, 836375400,
    836376300, 836377200, 836378100, 836379000, 836379900, 836380800,
    836381700, 836382600, 836383500, 836384400, 836385300, 836386200,
    836387100, 836388000, 836388900, 836389800, 836390700, 836391600,
    836392500, 836393400, 836394300, 836395200, 836396100, 836397000,
    836397900, 836398800, 836399700, 836400600, 836401500, 836402400,
    836403300, 836404200, 836405100, 836406000, 836406900, 836407800,
    836408700, 836409600, 836410500, 836411400, 836412300, 836413200,
    836414100, 836415000, 836415900, 836416800, 836417700, 836418600,
    836419500, 836420400, 836421300, 836422200, 836423100, 836424000,
    836424900, 836425800, 836426700, 836427600, 836428500, 836429400,
    836430300, 836431200, 836432100, 836433000, 836433900, 836434800,
    836435700, 836436600, 836437500, 836438400, 836439300, 836440200,
    836441100, 836442000, 836442900, 836443800, 836444700, 836445600,
    836446500, 836447400, 836448300, 836449200, 836450100, 836451000,
    836451900, 836452800, 836453700, 836454600, 836455500, 836456400,
    836457300, 836458200, 836459100, 836460000, 836460900, 836461800,
    836462700, 836463600, 836464500, 836465400, 836466300, 836467200,
    836468100, 836469000, 836469900, 836470800, 836471700, 836472600,
    836473500, 836474400, 836475300, 836476200, 836477100, 836478000,
    836478900, 836479800, 836480700, 836481600, 836482500, 836483400,
    836484300, 836485200, 836486100, 836487000, 836487900, 836488800,
    836489700, 836490600, 836491500, 836492400, 836493300, 836494200,
    836495100, 836496000, 836496900, 836497800, 836498700, 836499600,
    836500500, 836501400, 836502300, 836503200, 836504100, 836505000,
    836505900, 836506800, 836507700, 836508600, 836509500, 836510400,
    836511300, 836512200, 836513100, 836514000, 836514900, 836515800,
    836516700, 836517600, 836518500, 836519400, 836520300, 836521200,
    836522100, 836523000, 836523900, 836524800, 836525700, 836526600,
    836527500, 836528400, 836529300, 836530200, 836531100, 836532000,
    836532900, 836533800, 836534700, 836535600, 836536500, 836537400,
    836538300, 836539200, 836540100, 836541000, 836541900, 836542800,
    836543700, 836544600, 836545500, 836546400, 836547300, 836548200,
    836549100, 836550000, 836550900, 836551800, 836552700, 836553600,
    836554500, 836555400, 836556300, 836557200, 836558100, 836559000,
    836559900, 836560800, 836561700, 836562600, 836563500, 836564400,
    836565300, 836566200, 836567100, 836568000, 836568900, 836569800,
    836570700, 836571600, 836572500, 836573400, 836574300, 836575200,
    836576100, 836577000, 836577900, 836578800, 836579700, 836580600,
    836581500, 836582400, 836583300, 836584200, 836585100, 836586000,
    836586900, 836587800, 836588700, 836589600, 836590500, 836591400,
    836592300, 836593200, 836594100, 836595000, 836595900, 836596800,
    836597700, 836598600, 836599500, 836600400, 836601300, 836602200,
    836603100, 836604000, 836604900, 836605800, 836606700, 836607600,
    836608500, 836609400, 836610300, 836611200, 836612100, 836613000,
    836613900, 836614800, 836615700, 836616600, 836617500, 836618400,
    836619300, 836620200, 836621100, 836622000, 836622900, 836623800,
    836624700, 836625600, 836626500, 836627400, 836628300, 836629200,
    836630100, 836631000, 836631900, 836632800, 836633700, 836634600,
    836635500, 836636400, 836637300, 836638200, 836639100, 836640000,
    836640900, 836641800, 836642700, 836643600, 836644500, 836645400,
    836646300, 836647200, 836648100, 836649000, 836649900, 836650800,
    836651700, 836652600, 836653500, 836654400, 836655300, 836656200,
    836657100, 836658000, 836658900, 836659800, 836660700, 836661600,
    836662500, 836663400, 836664300, 836665200, 836666100, 836667000,
    836667900, 836668800, 836669700, 836670600, 836671500, 836672400,
    836673300, 836674200, 836675100, 836676000, 836676900, 836677800,
    836678700, 836679600, 836680500, 836681400, 836682300, 836683200,
    836684100, 836685000, 836685900, 836686800, 836687700, 836688600,
    836689500, 836690400, 836691300, 836692200, 836693100, 836694000,
    836694900, 836695800, 836696700, 836697600, 836698500, 836699400,
    836700300, 836701200, 836702100, 836703000, 836703900, 836704800,
    836705700, 836706600, 836707500, 836708400, 836709300, 836710200,
    836711100, 836712000, 836712900, 836713800, 836714700, 836715600,
    836716500, 836717400, 836718300, 836719200, 836720100, 836721000,
    836721900, 836722800, 836723700, 836724600, 836725500, 836726400,
    836727300, 836728200, 836729100, 836730000, 836730900, 836731800,
    836732700, 836733600, 836734500, 836735400, 836736300, 836737200,
    836738100, 836739000, 836739900, 836740800, 836741700, 836742600,
    836743500, 836744400, 836745300, 836746200, 836747100, 836748000,
    836748900, 836749800, 836750700, 836751600, 836752500, 836753400,
    836754300, 836755200, 836756100, 836757000, 836757900, 836758800,
    836759700, 836760600, 836761500, 836762400, 836763300, 836764200,
    836765100, 836766000, 836766900, 836767800, 836768700, 836769600,
    836770500, 836771400, 836772300, 836773200, 836774100, 836775000,
    836775900, 836776800, 836777700, 836778600, 836779500, 836780400,
    836781300, 836782200, 836783100, 836784000, 836784900, 836785800,
    836786700, 836787600, 836788500, 836789400, 836790300, 836791200,
    836792100, 836793000, 836793900, 836794800, 836795700, 836796600,
    836797500, 836798400, 836799300, 836800200, 836801100, 836802000,
    836802900, 836803800, 836804700, 836805600, 836806500, 836807400,
    836808300, 836809200, 836810100, 836811000, 836811900, 836812800,
    836813700, 836814600, 836815500, 836816400, 836817300, 836818200,
    836819100, 836820000, 836820900, 836821800, 836822700, 836823600,
    836824500, 836825400, 836826300, 836827200, 836828100, 836829000,
    836829900, 836830800, 836831700, 836832600, 836833500, 836834400,
    836835300, 836836200, 836837100, 836838000, 836838900, 836839800,
    836840700, 836841600, 836842500, 836843400, 836844300, 836845200,
    836846100, 836847000, 836847900, 836848800, 836849700, 836850600,
    836851500, 836852400, 836853300, 836854200, 836855100, 836856000,
    836856900, 836857800, 836858700, 836859600, 836860500, 836861400,
    836862300, 836863200, 836864100, 836865000, 836865900, 836866800,
    836867700, 836868600, 836869500, 836870400, 836871300, 836872200,
    836873100, 836874000, 836874900, 836875800, 836876700, 836877600,
    836878500, 836879400, 836880300, 836881200, 836882100, 836883000,
    836883900, 836884800, 836885700, 836886600, 836887500, 836888400,
    836889300, 836890200, 836891100, 836892000, 836892900, 836893800,
    836894700, 836895600, 836896500, 836897400, 836898300, 836899200,
    836900100, 836901000, 836901900, 836902800, 836903700, 836904600,
    836905500, 836906400, 836907300, 836908200, 836909100, 836910000,
    836910900, 836911800, 836912700, 836913600, 836914500, 836915400,
    836916300, 836917200, 836918100, 836919000, 836919900, 836920800,
    836921700, 836922600, 836923500, 836924400, 836925300, 836926200,
    836927100, 836928000, 836928900, 836929800, 836930700, 836931600,
    836932500, 836933400, 836934300, 836935200, 836936100, 836937000,
    836937900, 836938800, 836939700, 836940600, 836941500, 836942400,
    836943300, 836944200, 836945100, 836946000, 836946900, 836947800,
    836948700, 836949600, 836950500, 836951400, 836952300, 836953200,
    836954100, 836955000, 836955900, 836956800, 836957700, 836958600,
    836959500, 836960400, 836961300, 836962200, 836963100, 836964000,
    836964900, 836965800, 836966700, 836967600, 836968500, 836969400,
    836970300, 836971200, 836972100, 836973000, 836973900, 836974800,
    836975700, 836976600, 836977500, 836978400, 836979300, 836980200,
    836981100, 836982000, 836982900, 836983800, 836984700, 836985600,
    836986500, 836987400, 836988300, 836989200, 836990100, 836991000,
    836991900, 836992800, 836993700, 836994600, 836995500, 836996400,
    836997300, 836998200, 836999100, 837000000, 837000900, 837001800,
    837002700, 837003600, 837004500, 837005400, 837006300, 837007200,
    837008100, 837009000, 837009900, 837010800, 837011700, 837012600,
    837013500, 837014400, 837015300, 837016200, 837017100, 837018000,
    837018900, 837019800, 837020700, 837021600, 837022500, 837023400,
    837024300, 837025200, 837026100, 837027000, 837027900, 837028800,
    837029700, 837030600, 837031500, 837032400, 837033300, 837034200,
    837035100, 837036000, 837036900, 837037800, 837038700, 837039600,
    837040500, 837041400, 837042300, 837043200, 837044100, 837045000,
    837045900, 837046800, 837047700, 837048600, 837049500, 837050400,
    837051300, 837052200, 837053100, 837054000, 837054900, 837055800,
    837056700, 837057600, 837058500, 837059400, 837060300, 837061200,
    837062100, 837063000, 837063900, 837064800, 837065700, 837066600,
    837067500, 837068400, 837069300, 837070200, 837071100, 837072000,
    837072900, 837073800, 837074700, 837075600, 837076500, 837077400,
    837078300, 837079200, 837080100, 837081000, 837081900, 837082800,
    837083700, 837084600, 837085500, 837086400, 837087300, 837088200,
    837089100, 837090000, 837090900, 837091800, 837092700, 837093600,
    837094500, 837095400, 837096300, 837097200, 837098100, 837099000,
    837099900, 837100800, 837101700, 837102600, 837103500, 837104400,
    837105300, 837106200, 837107100, 837108000, 837108900, 837109800,
    837110700, 837111600, 837112500, 837113400, 837114300, 837115200,
    837116100, 837117000, 837117900, 837118800, 837119700, 837120600,
    837121500, 837122400, 837123300, 837124200, 837125100, 837126000,
    837126900, 837127800, 837128700, 837129600, 837130500, 837131400,
    837132300, 837133200, 837134100, 837135000, 837135900, 837136800,
    837137700, 837138600, 837139500, 837140400, 837141300, 837142200,
    837143100, 837144000, 837144900, 837145800, 837146700, 837147600,
    837148500, 837149400, 837150300, 837151200, 837152100, 837153000,
    837153900, 837154800, 837155700, 837156600, 837157500, 837158400,
    837159300, 837160200, 837161100, 837162000, 837162900, 837163800,
    837164700, 837165600, 837166500, 837167400, 837168300, 837169200,
    837170100, 837171000, 837171900, 837172800, 837173700, 837174600,
    837175500, 837176400, 837177300, 837178200, 837179100, 837180000,
    837180900, 837181800, 837182700, 837183600, 837184500, 837185400,
    837186300, 837187200, 837188100, 837189000, 837189900, 837190800,
    837191700, 837192600, 837193500, 837194400, 837195300, 837196200,
    837197100, 837198000, 837198900, 837199800, 837200700, 837201600,
    837202500, 837203400, 837204300, 837205200, 837206100, 837207000,
    837207900, 837208800, 837209700, 837210600, 837211500, 837212400,
    837213300, 837214200, 837215100, 837216000, 837216900, 837217800,
    837218700, 837219600, 837220500, 837221400, 837222300, 837223200,
    837224100, 837225000, 837225900, 837226800, 837227700, 837228600,
    837229500, 837230400, 837231300, 837232200, 837233100, 837234000,
    837234900, 837235800, 837236700, 837237600, 837238500, 837239400,
    837240300, 837241200, 837242100, 837243000, 837243900, 837244800,
    837245700, 837246600, 837247500, 837248400, 837249300, 837250200,
    837251100, 837252000, 837252900, 837253800, 837254700, 837255600,
    837256500, 837257400, 837258300, 837259200, 837260100, 837261000,
    837261900, 837262800, 837263700, 837264600, 837265500, 837266400,
    837267300, 837268200, 837269100, 837270000, 837270900, 837271800,
    837272700, 837273600, 837274500, 837275400, 837276300, 837277200,
    837278100, 837279000, 837279900, 837280800, 837281700, 837282600,
    837283500, 837284400, 837285300, 837286200, 837287100, 837288000,
    837288900, 837289800, 837290700, 837291600, 837292500, 837293400,
    837294300, 837295200, 837296100, 837297000, 837297900, 837298800,
    837299700, 837300600, 837301500, 837302400, 837303300, 837304200,
    837305100, 837306000, 837306900, 837307800, 837308700, 837309600,
    837310500, 837311400, 837312300, 837313200, 837314100, 837315000,
    837315900, 837316800, 837317700, 837318600, 837319500, 837320400,
    837321300, 837322200, 837323100, 837324000, 837324900, 837325800,
    837326700, 837327600, 837328500, 837329400, 837330300, 837331200,
    837332100, 837333000, 837333900, 837334800, 837335700, 837336600,
    837337500, 837338400, 837339300, 837340200, 837341100, 837342000,
    837342900, 837343800, 837344700, 837345600, 837346500, 837347400,
    837348300, 837349200, 837350100, 837351000, 837351900, 837352800,
    837353700, 837354600, 837355500, 837356400, 837357300, 837358200,
    837359100, 837360000, 837360900, 837361800, 837362700, 837363600,
    837364500, 837365400, 837366300, 837367200, 837368100, 837369000,
    837369900, 837370800, 837371700, 837372600, 837373500, 837374400,
    837375300, 837376200, 837377100, 837378000, 837378900, 837379800,
    837380700, 837381600, 837382500, 837383400, 837384300, 837385200,
    837386100, 837387000, 837387900, 837388800, 837389700, 837390600,
    837391500, 837392400, 837393300, 837394200, 837395100, 837396000,
    837396900, 837397800, 837398700, 837399600, 837400500, 837401400,
    837402300, 837403200, 837404100, 837405000, 837405900, 837406800,
    837407700, 837408600, 837409500, 837410400, 837411300, 837412200,
    837413100, 837414000, 837414900, 837415800, 837416700, 837417600,
    837418500, 837419400, 837420300, 837421200, 837422100, 837423000,
    837423900, 837424800, 837425700, 837426600, 837427500, 837428400,
    837429300, 837430200, 837431100, 837432000, 837432900, 837433800,
    837434700, 837435600, 837436500, 837437400, 837438300, 837439200,
    837440100, 837441000, 837441900, 837442800, 837443700, 837444600,
    837445500, 837446400, 837447300, 837448200, 837449100, 837450000,
    837450900, 837451800, 837452700, 837453600, 837454500, 837455400,
    837456300, 837457200, 837458100, 837459000, 837459900, 837460800,
    837461700, 837462600, 837463500, 837464400, 837465300, 837466200,
    837467100, 837468000, 837468900, 837469800, 837470700, 837471600,
    837472500, 837473400, 837474300, 837475200, 837476100, 837477000,
    837477900, 837478800, 837479700, 837480600, 837481500, 837482400,
    837483300, 837484200, 837485100, 837486000, 837486900, 837487800,
    837488700, 837489600, 837490500, 837491400, 837492300, 837493200,
    837494100, 837495000, 837495900, 837496800, 837497700, 837498600,
    837499500, 837500400, 837501300, 837502200, 837503100, 837504000,
    837504900, 837505800, 837506700, 837507600, 837508500, 837509400,
    837510300, 837511200, 837512100, 837513000, 837513900, 837514800,
    837515700, 837516600, 837517500, 837518400, 837519300, 837520200,
    837521100, 837522000, 837522900, 837523800, 837524700, 837525600,
    837526500, 837527400, 837528300, 837529200, 837530100, 837531000,
    837531900, 837532800, 837533700, 837534600, 837535500, 837536400,
    837537300, 837538200, 837539100, 837540000, 837540900, 837541800,
    837542700, 837543600, 837544500, 837545400, 837546300, 837547200,
    837548100, 837549000, 837549900, 837550800, 837551700, 837552600,
    837553500, 837554400, 837555300, 837556200, 837557100, 837558000,
    837558900, 837559800, 837560700, 837561600, 837562500, 837563400,
    837564300, 837565200, 837566100, 837567000, 837567900, 837568800,
    837569700, 837570600, 837571500, 837572400, 837573300, 837574200,
    837575100, 837576000, 837576900, 837577800, 837578700, 837579600,
    837580500, 837581400, 837582300, 837583200, 837584100, 837585000,
    837585900, 837586800, 837587700, 837588600, 837589500, 837590400,
    837591300, 837592200, 837593100, 837594000, 837594900, 837595800,
    837596700, 837597600, 837598500, 837599400, 837600300, 837601200,
    837602100, 837603000, 837603900, 837604800, 837605700, 837606600,
    837607500, 837608400, 837609300, 837610200, 837611100, 837612000,
    837612900, 837613800, 837614700, 837615600, 837616500, 837617400,
    837618300, 837619200, 837620100, 837621000, 837621900, 837622800,
    837623700, 837624600, 837625500, 837626400, 837627300, 837628200,
    837629100, 837630000, 837630900, 837631800, 837632700, 837633600,
    837634500, 837635400, 837636300, 837637200, 837638100, 837639000,
    837639900, 837640800, 837641700, 837642600, 837643500, 837644400,
    837645300, 837646200, 837647100, 837648000, 837648900, 837649800,
    837650700, 837651600, 837652500, 837653400, 837654300, 837655200,
    837656100, 837657000, 837657900, 837658800, 837659700, 837660600,
    837661500, 837662400, 837663300, 837664200, 837665100, 837666000,
    837666900, 837667800, 837668700, 837669600, 837670500, 837671400,
    837672300, 837673200, 837674100, 837675000, 837675900, 837676800,
    837677700, 837678600, 837679500, 837680400, 837681300, 837682200,
    837683100, 837684000, 837684900, 837685800, 837686700, 837687600,
    837688500, 837689400, 837690300, 837691200, 837692100, 837693000,
    837693900, 837694800, 837695700, 837696600, 837697500, 837698400,
    837699300, 837700200, 837701100, 837702000, 837702900, 837703800,
    837704700, 837705600, 837706500, 837707400, 837708300, 837709200,
    837710100, 837711000, 837711900, 837712800, 837713700, 837714600,
    837715500, 837716400, 837717300, 837718200, 837719100, 837720000,
    837720900, 837721800, 837722700, 837723600, 837724500, 837725400,
    837726300, 837727200, 837728100, 837729000, 837729900, 837730800,
    837731700, 837732600, 837733500, 837734400, 837735300, 837736200,
    837737100, 837738000, 837738900, 837739800, 837740700, 837741600,
    837742500, 837743400, 837744300, 837745200, 837746100, 837747000,
    837747900, 837748800, 837749700, 837750600, 837751500, 837752400,
    837753300, 837754200, 837755100, 837756000, 837756900, 837757800,
    837758700, 837759600, 837760500, 837761400, 837762300, 837763200,
    837764100, 837765000, 837765900, 837766800, 837767700, 837768600,
    837769500, 837770400, 837771300, 837772200, 837773100, 837774000,
    837774900, 837775800, 837776700, 837777600, 837778500, 837779400,
    837780300, 837781200, 837782100, 837783000, 837783900, 837784800,
    837785700, 837786600, 837787500, 837788400, 837789300, 837790200,
    837791100, 837792000, 837792900, 837793800, 837794700, 837795600,
    837796500, 837797400, 837798300, 837799200, 837800100, 837801000,
    837801900, 837802800, 837803700, 837804600, 837805500, 837806400,
    837807300, 837808200, 837809100, 837810000, 837810900, 837811800,
    837812700, 837813600, 837814500, 837815400, 837816300, 837817200,
    837818100, 837819000, 837819900, 837820800, 837821700, 837822600,
    837823500, 837824400, 837825300, 837826200, 837827100, 837828000,
    837828900, 837829800, 837830700, 837831600, 837832500, 837833400,
    837834300, 837835200, 837836100, 837837000, 837837900, 837838800,
    837839700, 837840600, 837841500, 837842400, 837843300, 837844200,
    837845100, 837846000, 837846900, 837847800, 837848700, 837849600,
    837850500, 837851400, 837852300, 837853200, 837854100, 837855000,
    837855900, 837856800, 837857700, 837858600, 837859500, 837860400,
    837861300, 837862200, 837863100, 837864000, 837864900, 837865800,
    837866700, 837867600, 837868500, 837869400, 837870300, 837871200,
    837872100, 837873000, 837873900, 837874800, 837875700, 837876600,
    837877500, 837878400, 837879300, 837880200, 837881100, 837882000,
    837882900, 837883800, 837884700, 837885600, 837886500, 837887400,
    837888300, 837889200, 837890100, 837891000, 837891900, 837892800,
    837893700, 837894600, 837895500, 837896400, 837897300, 837898200,
    837899100, 837900000, 837900900, 837901800, 837902700, 837903600,
    837904500, 837905400, 837906300, 837907200, 837908100, 837909000,
    837909900, 837910800, 837911700, 837912600, 837913500, 837914400,
    837915300, 837916200, 837917100, 837918000, 837918900, 837919800,
    837920700, 837921600, 837922500, 837923400, 837924300, 837925200,
    837926100, 837927000, 837927900, 837928800, 837929700, 837930600,
    837931500, 837932400, 837933300, 837934200, 837935100, 837936000,
    837936900, 837937800, 837938700, 837939600, 837940500, 837941400,
    837942300, 837943200, 837944100, 837945000, 837945900, 837946800,
    837947700, 837948600, 837949500, 837950400, 837951300, 837952200,
    837953100, 837954000, 837954900, 837955800, 837956700, 837957600,
    837958500, 837959400, 837960300, 837961200, 837962100, 837963000,
    837963900, 837964800, 837965700, 837966600, 837967500, 837968400,
    837969300, 837970200, 837971100, 837972000, 837972900, 837973800,
    837974700, 837975600, 837976500, 837977400, 837978300, 837979200,
    837980100, 837981000, 837981900, 837982800, 837983700, 837984600,
    837985500, 837986400, 837987300, 837988200, 837989100, 837990000,
    837990900, 837991800, 837992700, 837993600, 837994500, 837995400,
    837996300, 837997200, 837998100, 837999000, 837999900, 838000800,
    838001700, 838002600, 838003500, 838004400, 838005300, 838006200,
    838007100, 838008000, 838008900, 838009800, 838010700, 838011600,
    838012500, 838013400, 838014300, 838015200, 838016100, 838017000,
    838017900, 838018800, 838019700, 838020600, 838021500, 838022400,
    838023300, 838024200, 838025100, 838026000, 838026900, 838027800,
    838028700, 838029600, 838030500, 838031400, 838032300, 838033200,
    838034100, 838035000, 838035900, 838036800, 838037700, 838038600,
    838039500, 838040400, 838041300, 838042200, 838043100, 838044000,
    838044900, 838045800, 838046700, 838047600, 838048500, 838049400,
    838050300, 838051200, 838052100, 838053000, 838053900, 838054800,
    838055700, 838056600, 838057500, 838058400, 838059300, 838060200,
    838061100, 838062000, 838062900, 838063800, 838064700, 838065600,
    838066500, 838067400, 838068300, 838069200, 838070100, 838071000,
    838071900, 838072800, 838073700, 838074600, 838075500, 838076400,
    838077300, 838078200, 838079100, 838080000, 838080900, 838081800,
    838082700, 838083600, 838084500, 838085400, 838086300, 838087200,
    838088100, 838089000, 838089900, 838090800, 838091700, 838092600,
    838093500, 838094400, 838095300, 838096200, 838097100, 838098000,
    838098900, 838099800, 838100700, 838101600, 838102500, 838103400,
    838104300, 838105200, 838106100, 838107000, 838107900, 838108800,
    838109700, 838110600, 838111500, 838112400, 838113300, 838114200,
    838115100, 838116000, 838116900, 838117800, 838118700, 838119600,
    838120500, 838121400, 838122300, 838123200, 838124100, 838125000,
    838125900, 838126800, 838127700, 838128600, 838129500, 838130400,
    838131300, 838132200, 838133100, 838134000, 838134900, 838135800,
    838136700, 838137600, 838138500, 838139400, 838140300, 838141200,
    838142100, 838143000, 838143900, 838144800, 838145700, 838146600,
    838147500, 838148400, 838149300, 838150200, 838151100, 838152000,
    838152900, 838153800, 838154700, 838155600, 838156500, 838157400,
    838158300, 838159200, 838160100, 838161000, 838161900, 838162800,
    838163700, 838164600, 838165500, 838166400, 838167300, 838168200,
    838169100, 838170000, 838170900, 838171800, 838172700, 838173600,
    838174500, 838175400, 838176300, 838177200, 838178100, 838179000,
    838179900, 838180800, 838181700, 838182600, 838183500, 838184400,
    838185300, 838186200, 838187100, 838188000, 838188900, 838189800,
    838190700, 838191600, 838192500, 838193400, 838194300, 838195200,
    838196100, 838197000, 838197900, 838198800, 838199700, 838200600,
    838201500, 838202400, 838203300, 838204200, 838205100, 838206000,
    838206900, 838207800, 838208700, 838209600, 838210500, 838211400,
    838212300, 838213200, 838214100, 838215000, 838215900, 838216800,
    838217700, 838218600, 838219500, 838220400, 838221300, 838222200,
    838223100, 838224000, 838224900, 838225800, 838226700, 838227600,
    838228500, 838229400, 838230300, 838231200, 838232100, 838233000,
    838233900, 838234800, 838235700, 838236600, 838237500, 838238400,
    838239300, 838240200, 838241100, 838242000, 838242900, 838243800,
    838244700, 838245600, 838246500, 838247400, 838248300, 838249200,
    838250100, 838251000, 838251900, 838252800, 838253700, 838254600,
    838255500, 838256400, 838257300, 838258200, 838259100, 838260000,
    838260900, 838261800, 838262700, 838263600, 838264500, 838265400,
    838266300, 838267200, 838268100, 838269000, 838269900, 838270800,
    838271700, 838272600, 838273500, 838274400, 838275300, 838276200,
    838277100, 838278000, 838278900, 838279800, 838280700, 838281600,
    838282500, 838283400, 838284300, 838285200, 838286100, 838287000,
    838287900, 838288800, 838289700, 838290600, 838291500, 838292400,
    838293300, 838294200, 838295100, 838296000, 838296900, 838297800,
    838298700, 838299600, 838300500, 838301400, 838302300, 838303200,
    838304100, 838305000, 838305900, 838306800, 838307700, 838308600,
    838309500, 838310400, 838311300, 838312200, 838313100, 838314000,
    838314900, 838315800, 838316700, 838317600, 838318500, 838319400,
    838320300, 838321200, 838322100, 838323000, 838323900, 838324800,
    838325700, 838326600, 838327500, 838328400, 838329300, 838330200,
    838331100, 838332000, 838332900, 838333800, 838334700, 838335600,
    838336500, 838337400, 838338300, 838339200, 838340100, 838341000,
    838341900, 838342800, 838343700, 838344600, 838345500, 838346400,
    838347300, 838348200, 838349100, 838350000, 838350900, 838351800,
    838352700, 838353600, 838354500, 838355400, 838356300, 838357200,
    838358100, 838359000, 838359900, 838360800, 838361700, 838362600,
    838363500, 838364400, 838365300, 838366200, 838367100, 838368000,
    838368900, 838369800, 838370700, 838371600, 838372500, 838373400,
    838374300, 838375200, 838376100, 838377000, 838377900, 838378800,
    838379700, 838380600, 838381500, 838382400, 838383300, 838384200,
    838385100, 838386000, 838386900, 838387800, 838388700, 838389600,
    838390500, 838391400, 838392300, 838393200, 838394100, 838395000,
    838395900, 838396800, 838397700, 838398600, 838399500, 838400400,
    838401300, 838402200, 838403100, 838404000, 838404900, 838405800,
    838406700, 838407600, 838408500, 838409400, 838410300, 838411200,
    838412100, 838413000, 838413900, 838414800, 838415700, 838416600,
    838417500, 838418400, 838419300, 838420200, 838421100, 838422000,
    838422900, 838423800, 838424700, 838425600, 838426500, 838427400,
    838428300, 838429200, 838430100, 838431000, 838431900, 838432800,
    838433700, 838434600, 838435500, 838436400, 838437300, 838438200,
    838439100, 838440000, 838440900, 838441800, 838442700, 838443600,
    838444500, 838445400, 838446300, 838447200, 838448100, 838449000,
    838449900, 838450800, 838451700, 838452600, 838453500, 838454400,
    838455300, 838456200, 838457100, 838458000, 838458900, 838459800,
    838460700, 838461600, 838462500, 838463400, 838464300, 838465200,
    838466100, 838467000, 838467900, 838468800, 838469700, 838470600,
    838471500, 838472400, 838473300, 838474200, 838475100, 838476000,
    838476900, 838477800, 838478700, 838479600, 838480500, 838481400,
    838482300, 838483200, 838484100, 838485000, 838485900, 838486800,
    838487700, 838488600, 838489500, 838490400, 838491300, 838492200,
    838493100, 838494000, 838494900, 838495800, 838496700, 838497600,
    838498500, 838499400, 838500300, 838501200, 838502100, 838503000,
    838503900, 838504800, 838505700, 838506600, 838507500, 838508400,
    838509300, 838510200, 838511100, 838512000, 838512900, 838513800,
    838514700, 838515600, 838516500, 838517400, 838518300, 838519200,
    838520100, 838521000, 838521900, 838522800, 838523700, 838524600,
    838525500, 838526400, 838527300, 838528200, 838529100, 838530000,
    838530900, 838531800, 838532700, 838533600, 838534500, 838535400,
    838536300, 838537200, 838538100, 838539000, 838539900, 838540800,
    838541700, 838542600, 838543500, 838544400, 838545300, 838546200,
    838547100, 838548000, 838548900, 838549800, 838550700, 838551600,
    838552500, 838553400, 838554300, 838555200, 838556100, 838557000,
    838557900, 838558800, 838559700, 838560600, 838561500, 838562400,
    838563300, 838564200, 838565100, 838566000, 838566900, 838567800,
    838568700, 838569600, 838570500, 838571400, 838572300, 838573200,
    838574100, 838575000, 838575900, 838576800, 838577700, 838578600,
    838579500, 838580400, 838581300, 838582200, 838583100, 838584000,
    838584900, 838585800, 838586700, 838587600, 838588500, 838589400,
    838590300, 838591200, 838592100, 838593000, 838593900, 838594800,
    838595700, 838596600, 838597500, 838598400, 838599300, 838600200,
    838601100, 838602000, 838602900, 838603800, 838604700, 838605600,
    838606500, 838607400, 838608300, 838609200, 838610100, 838611000,
    838611900, 838612800, 838613700, 838614600, 838615500, 838616400,
    838617300, 838618200, 838619100, 838620000, 838620900, 838621800,
    838622700, 838623600, 838624500, 838625400, 838626300, 838627200,
    838628100, 838629000, 838629900, 838630800, 838631700, 838632600,
    838633500, 838634400, 838635300, 838636200, 838637100, 838638000,
    838638900, 838639800, 838640700, 838641600, 838642500, 838643400,
    838644300, 838645200, 838646100, 838647000, 838647900, 838648800,
    838649700, 838650600, 838651500, 838652400, 838653300, 838654200,
    838655100, 838656000, 838656900, 838657800, 838658700, 838659600,
    838660500, 838661400, 838662300, 838663200, 838664100, 838665000,
    838665900, 838666800, 838667700, 838668600, 838669500, 838670400,
    838671300, 838672200, 838673100, 838674000, 838674900, 838675800,
    838676700, 838677600, 838678500, 838679400, 838680300, 838681200,
    838682100, 838683000, 838683900, 838684800, 838685700, 838686600,
    838687500, 838688400, 838689300, 838690200, 838691100, 838692000,
    838692900, 838693800, 838694700, 838695600, 838696500, 838697400,
    838698300, 838699200, 838700100, 838701000, 838701900, 838702800,
    838703700, 838704600, 838705500, 838706400, 838707300, 838708200,
    838709100, 838710000, 838710900, 838711800, 838712700, 838713600,
    838714500, 838715400, 838716300, 838717200, 838718100, 838719000,
    838719900, 838720800, 838721700, 838722600, 838723500, 838724400,
    838725300, 838726200, 838727100, 838728000, 838728900, 838729800,
    838730700, 838731600, 838732500, 838733400, 838734300, 838735200,
    838736100, 838737000, 838737900, 838738800, 838739700, 838740600,
    838741500, 838742400, 838743300, 838744200, 838745100, 838746000,
    838746900, 838747800, 838748700, 838749600, 838750500, 838751400,
    838752300, 838753200, 838754100, 838755000, 838755900, 838756800,
    838757700, 838758600, 838759500, 838760400, 838761300, 838762200,
    838763100, 838764000, 838764900, 838765800, 838766700, 838767600,
    838768500, 838769400, 838770300, 838771200, 838772100, 838773000,
    838773900, 838774800, 838775700, 838776600, 838777500, 838778400,
    838779300, 838780200, 838781100, 838782000, 838782900, 838783800,
    838784700, 838785600, 838786500, 838787400, 838788300, 838789200,
    838790100, 838791000, 838791900, 838792800, 838793700, 838794600,
    838795500, 838796400, 838797300, 838798200, 838799100, 838800000,
    838800900, 838801800, 838802700, 838803600, 838804500, 838805400,
    838806300, 838807200, 838808100, 838809000, 838809900, 838810800,
    838811700, 838812600, 838813500, 838814400, 838815300, 838816200,
    838817100, 838818000, 838818900, 838819800, 838820700, 838821600,
    838822500, 838823400, 838824300, 838825200, 838826100, 838827000,
    838827900, 838828800, 838829700, 838830600, 838831500, 838832400,
    838833300, 838834200, 838835100, 838836000, 838836900, 838837800,
    838838700, 838839600, 838840500, 838841400, 838842300, 838843200,
    838844100, 838845000, 838845900, 838846800, 838847700, 838848600,
    838849500, 838850400, 838851300, 838852200, 838853100, 838854000,
    838854900, 838855800, 838856700, 838857600, 838858500, 838859400,
    838860300, 838861200, 838862100, 838863000, 838863900, 838864800,
    838865700, 838866600, 838867500, 838868400, 838869300, 838870200,
    838871100, 838872000, 838872900, 838873800, 838874700, 838875600,
    838876500, 838877400, 838878300, 838879200, 838880100, 838881000,
    838881900, 838882800, 838883700, 838884600, 838885500, 838886400,
    838887300, 838888200, 838889100, 838890000, 838890900, 838891800,
    838892700, 838893600, 838894500, 838895400, 838896300, 838897200,
    838898100, 838899000, 838899900, 838900800, 838901700, 838902600,
    838903500, 838904400, 838905300, 838906200, 838907100, 838908000,
    838908900, 838909800, 838910700, 838911600, 838912500, 838913400,
    838914300, 838915200, 838916100, 838917000, 838917900, 838918800,
    838919700, 838920600, 838921500, 838922400, 838923300, 838924200,
    838925100, 838926000, 838926900, 838927800, 838928700, 838929600,
    838930500, 838931400, 838932300, 838933200, 838934100, 838935000,
    838935900, 838936800, 838937700, 838938600, 838939500, 838940400,
    838941300, 838942200, 838943100, 838944000, 838944900, 838945800,
    838946700, 838947600, 838948500, 838949400, 838950300, 838951200,
    838952100, 838953000, 838953900, 838954800, 838955700, 838956600,
    838957500, 838958400, 838959300, 838960200, 838961100, 838962000,
    838962900, 838963800, 838964700, 838965600, 838966500, 838967400,
    838968300, 838969200, 838970100, 838971000, 838971900, 838972800,
    838973700, 838974600, 838975500, 838976400, 838977300, 838978200,
    838979100, 838980000, 838980900, 838981800, 838982700, 838983600,
    838984500, 838985400, 838986300, 838987200, 838988100, 838989000,
    838989900, 838990800, 838991700, 838992600, 838993500, 838994400,
    838995300, 838996200, 838997100, 838998000, 838998900, 838999800,
    839000700, 839001600, 839002500, 839003400, 839004300, 839005200,
    839006100, 839007000, 839007900, 839008800, 839009700, 839010600,
    839011500, 839012400, 839013300, 839014200, 839015100, 839016000,
    839016900, 839017800, 839018700, 839019600, 839020500, 839021400,
    839022300, 839023200, 839024100, 839025000, 839025900, 839026800,
    839027700, 839028600, 839029500, 839030400, 839031300, 839032200,
    839033100, 839034000, 839034900, 839035800, 839036700, 839037600,
    839038500, 839039400, 839040300, 839041200, 839042100, 839043000,
    839043900, 839044800, 839045700, 839046600, 839047500, 839048400,
    839049300, 839050200, 839051100, 839052000, 839052900, 839053800,
    839054700, 839055600, 839056500, 839057400, 839058300, 839059200,
    839060100, 839061000, 839061900, 839062800, 839063700, 839064600,
    839065500, 839066400, 839067300, 839068200, 839069100, 839070000,
    839070900, 839071800, 839072700, 839073600, 839074500, 839075400,
    839076300, 839077200, 839078100, 839079000, 839079900, 839080800,
    839081700, 839082600, 839083500, 839084400, 839085300, 839086200,
    839087100, 839088000, 839088900, 839089800, 839090700, 839091600,
    839092500, 839093400, 839094300, 839095200, 839096100, 839097000,
    839097900, 839098800, 839099700, 839100600, 839101500, 839102400,
    839103300, 839104200, 839105100, 839106000, 839106900, 839107800,
    839108700, 839109600, 839110500, 839111400, 839112300, 839113200,
    839114100, 839115000, 839115900, 839116800, 839117700, 839118600,
    839119500, 839120400, 839121300, 839122200, 839123100, 839124000,
    839124900, 839125800, 839126700, 839127600, 839128500, 839129400,
    839130300, 839131200, 839132100, 839133000, 839133900, 839134800,
    839135700, 839136600, 839137500, 839138400, 839139300, 839140200,
    839141100, 839142000, 839142900, 839143800, 839144700, 839145600,
    839146500, 839147400, 839148300, 839149200, 839150100, 839151000,
    839151900, 839152800, 839153700, 839154600, 839155500, 839156400,
    839157300, 839158200, 839159100, 839160000, 839160900, 839161800,
    839162700, 839163600, 839164500, 839165400, 839166300, 839167200,
    839168100, 839169000, 839169900, 839170800, 839171700, 839172600,
    839173500, 839174400, 839175300, 839176200, 839177100, 839178000,
    839178900, 839179800, 839180700, 839181600, 839184300, 839185200,
    839186100, 839187000, 839187900, 839188800, 839189700, 839190600,
    839191500, 839192400, 839193300, 839194200, 839195100, 839196000,
    839196900, 839197800, 839198700, 839199600, 839200500, 839201400,
    839202300, 839203200, 839204100, 839205000, 839205900, 839206800,
    839207700, 839208600, 839209500, 839210400, 839211300, 839212200,
    839213100, 839214000, 839214900, 839215800, 839216700, 839217600,
    839218500, 839219400, 839220300, 839221200, 839222100, 839223000,
    839223900, 839224800, 839225700, 839226600, 839227500, 839228400,
    839229300, 839230200, 839231100, 839232000, 839232900, 839233800,
    839234700, 839235600, 839236500, 839237400, 839238300, 839239200,
    839240100, 839241000, 839241900, 839242800, 839243700, 839244600,
    839245500, 839246400, 839247300, 839248200, 839249100, 839250000,
    839250900, 839251800, 839252700, 839253600, 839254500, 839255400,
    839256300, 839257200, 839258100, 839259000, 839259900, 839260800,
    839261700, 839262600, 839263500, 839264400, 839265300, 839266200,
    839267100, 839268000, 839268900, 839269800, 839270700, 839271600,
    839272500, 839273400, 839274300, 839275200, 839276100, 839277000,
    839277900, 839278800, 839279700, 839280600, 839281500, 839282400,
    839283300, 839284200, 839285100, 839286000, 839286900, 839287800,
    839288700, 839289600, 839290500, 839291400, 839292300, 839293200,
    839294100, 839295000, 839295900, 839296800, 839297700, 839298600,
    839299500, 839300400, 839301300, 839302200, 839303100, 839304000,
    839304900, 839305800, 839306700, 839307600, 839308500, 839309400,
    839310300, 839311200, 839312100, 839313000, 839313900, 839314800,
    839315700, 839316600, 839317500, 839318400, 839319300, 839320200,
    839321100, 839322000, 839322900, 839323800, 839324700, 839325600,
    839326500, 839327400, 839328300, 839329200, 839330100, 839331000,
    839331900, 839332800, 839333700, 839334600, 839335500, 839336400,
    839337300, 839338200, 839339100, 839340000, 839340900, 839341800,
    839342700, 839343600, 839344500, 839345400, 839346300, 839347200,
    839348100, 839349000, 839349900, 839350800, 839351700, 839352600,
    839353500, 839354400, 839355300, 839356200, 839357100, 839358000,
    839358900, 839359800, 839360700, 839361600, 839362500, 839363400,
    839364300, 839365200, 839366100, 839367000, 839367900, 839368800,
    839369700, 839370600, 839371500, 839372400, 839373300, 839374200,
    839375100, 839376000, 839376900, 839377800, 839378700, 839379600,
    839380500, 839381400, 839382300, 839383200, 839384100, 839385000,
    839385900, 839386800, 839387700, 839388600, 839389500, 839390400,
    839391300, 839392200, 839393100, 839394000, 839394900, 839395800,
    839396700, 839397600, 839398500, 839399400, 839400300, 839401200,
    839402100, 839403000, 839403900, 839404800, 839405700, 839406600,
    839407500, 839408400, 839409300, 839410200, 839411100, 839412000,
    839412900, 839413800, 839414700, 839415600, 839416500, 839417400,
    839418300, 839419200, 839420100, 839421000, 839421900, 839422800,
    839423700, 839424600, 839425500, 839426400, 839427300, 839428200,
    839429100, 839430000, 839430900, 839431800, 839432700, 839433600,
    839434500, 839435400, 839436300, 839437200, 839438100, 839439000,
    839439900, 839440800, 839441700, 839442600, 839443500, 839444400,
    839445300, 839446200, 839447100, 839448000, 839448900, 839449800,
    839450700, 839451600, 839452500, 839453400, 839454300, 839455200,
    839456100, 839457000, 839457900, 839458800, 839459700, 839460600,
    839461500, 839462400, 839463300, 839464200, 839465100, 839466000,
    839466900, 839467800, 839468700, 839469600, 839470500, 839471400,
    839472300, 839473200, 839474100, 839475000, 839475900, 839476800,
    839477700, 839478600, 839479500, 839480400, 839481300, 839482200,
    839483100, 839484000, 839484900, 839485800, 839486700, 839487600,
    839488500, 839489400, 839490300, 839491200, 839492100, 839493000,
    839493900, 839494800, 839495700, 839496600, 839497500, 839498400,
    839499300, 839500200, 839501100, 839502000, 839502900, 839503800,
    839504700, 839505600, 839506500, 839507400, 839508300, 839509200,
    839510100, 839511000, 839511900, 839512800, 839513700, 839514600,
    839515500, 839516400, 839517300, 839518200, 839519100, 839520000,
    839520900, 839521800, 839522700, 839523600, 839524500, 839525400,
    839526300, 839527200, 839528100, 839529000, 839529900, 839530800,
    839531700, 839532600, 839533500, 839534400, 839535300, 839536200,
    839537100, 839538000, 839538900, 839539800, 839540700, 839541600,
    839542500, 839543400, 839544300, 839545200, 839546100, 839547000,
    839547900, 839548800, 839549700, 839550600, 839551500, 839552400,
    839553300, 839554200, 839555100, 839556000, 839556900, 839557800,
    839558700, 839559600, 839560500, 839561400, 839562300, 839563200,
    839564100, 839565000, 839565900, 839566800, 839567700, 839568600,
    839569500, 839570400, 839571300, 839572200, 839573100, 839574000,
    839574900, 839575800, 839576700, 839577600, 839578500, 839579400,
    839580300, 839581200, 839582100, 839583000, 839583900, 839584800,
    839585700, 839586600, 839587500, 839588400, 839589300, 839590200,
    839591100, 839592000, 839592900, 839593800, 839594700, 839595600,
    839596500, 839597400, 839598300, 839599200, 839600100, 839601000,
    839601900, 839602800, 839603700, 839604600, 839605500, 839606400,
    839607300, 839608200, 839609100, 839610000, 839610900, 839611800,
    839612700, 839613600, 839614500, 839615400, 839616300, 839617200,
    839618100, 839619000, 839619900, 839620800, 839621700, 839622600,
    839623500, 839624400, 839625300, 839626200, 839627100, 839628000,
    839628900, 839629800, 839630700, 839631600, 839632500, 839633400,
    839634300, 839635200, 839636100, 839637000, 839637900, 839638800,
    839639700, 839640600, 839641500, 839642400, 839643300, 839644200,
    839645100, 839646000, 839646900, 839647800, 839648700, 839649600,
    839650500, 839651400, 839652300, 839653200, 839654100, 839655000,
    839655900, 839656800, 839657700, 839658600, 839659500, 839660400,
    839661300, 839662200, 839663100, 839664000, 839664900, 839665800,
    839666700, 839667600, 839668500, 839669400, 839670300, 839671200,
    839672100, 839673000, 839673900, 839674800, 839675700, 839676600,
    839677500, 839678400, 839679300, 839680200, 839681100, 839682000,
    839682900, 839683800, 839684700, 839685600, 839686500, 839687400,
    839688300, 839689200, 839690100, 839691000, 839691900, 839692800,
    839693700, 839694600, 839695500, 839696400, 839697300, 839698200,
    839699100, 839700000, 839700900, 839701800, 839702700, 839703600,
    839704500, 839705400, 839706300, 839707200, 839708100, 839709000,
    839709900, 839710800, 839711700, 839712600, 839713500, 839714400,
    839715300, 839716200, 839717100, 839718000, 839718900, 839719800,
    839720700, 839721600, 839722500, 839723400, 839724300, 839725200,
    839726100, 839727000, 839727900, 839728800, 839729700, 839730600,
    839731500, 839732400, 839733300, 839734200, 839735100, 839736000,
    839736900, 839737800, 839738700, 839739600, 839740500, 839741400,
    839742300, 839743200, 839744100, 839745000, 839745900, 839746800,
    839747700, 839748600, 839749500, 839750400, 839751300, 839752200,
    839753100, 839754000, 839754900, 839755800, 839756700, 839757600,
    839758500, 839759400, 839760300, 839761200, 839762100, 839763000,
    839763900, 839764800, 839765700, 839766600, 839767500, 839768400,
    839769300, 839770200, 839771100, 839772000, 839772900, 839773800,
    839774700, 839775600, 839776500, 839777400, 839778300, 839779200,
    839780100, 839781000, 839781900, 839782800, 839783700, 839784600,
    839785500, 839786400, 839787300, 839788200, 839789100, 839790000,
    839790900, 839791800, 839792700, 839793600, 839794500, 839795400,
    839796300, 839797200, 839798100, 839799000, 839799900, 839800800,
    839801700, 839802600, 839803500, 839804400, 839805300, 839806200,
    839807100, 839808000, 839808900, 839809800, 839810700, 839811600,
    839812500, 839813400, 839814300, 839815200, 839816100, 839817000,
    839817900, 839818800, 839819700, 839820600, 839821500, 839822400,
    839823300, 839824200, 839825100, 839826000, 839826900, 839827800,
    839828700, 839829600, 839830500, 839831400, 839832300, 839833200,
    839834100, 839835000, 839835900, 839836800, 839837700, 839838600,
    839839500, 839840400, 839841300, 839842200, 839843100, 839844000,
    839844900, 839845800, 839846700, 839847600, 839848500, 839849400,
    839850300, 839851200, 839852100, 839853000, 839853900, 839854800,
    839855700, 839856600, 839857500, 839858400, 839859300, 839860200,
    839861100, 839862000, 839862900, 839863800, 839864700, 839865600,
    839866500, 839867400, 839868300, 839869200, 839870100, 839871000,
    839871900, 839872800, 839873700, 839874600, 839875500, 839876400,
    839877300, 839878200, 839879100, 839880000, 839880900, 839881800,
    839882700, 839883600, 839884500, 839885400, 839886300, 839887200,
    839888100, 839889000, 839889900, 839890800, 839891700, 839892600,
    839893500, 839894400, 839895300, 839896200, 839897100, 839898000,
    839898900, 839899800, 839900700, 839901600, 839902500, 839903400,
    839904300, 839905200, 839906100, 839907000, 839907900, 839908800,
    839909700, 839910600, 839911500, 839912400, 839913300, 839914200,
    839915100, 839916000, 839916900, 839917800, 839918700, 839919600,
    839920500, 839921400, 839922300, 839923200, 839924100, 839925000,
    839925900, 839926800, 839927700, 839928600, 839929500, 839930400,
    839931300, 839932200, 839933100, 839934000, 839934900, 839935800,
    839936700, 839937600, 839938500, 839939400, 839940300, 839941200,
    839942100, 839943000, 839943900, 839944800, 839945700, 839946600,
    839947500, 839948400, 839949300, 839950200, 839951100, 839952000,
    839952900, 839953800, 839954700, 839955600, 839956500, 839957400,
    839958300, 839959200, 839960100, 839961000, 839961900, 839962800,
    839963700, 839964600, 839965500, 839966400, 839967300, 839968200,
    839969100, 839970000, 839970900, 839971800, 839972700, 839973600,
    839974500, 839975400, 839976300, 839977200, 839978100, 839979000,
    839979900, 839980800, 839981700, 839982600, 839983500, 839984400,
    839985300, 839986200, 839987100, 839988000, 839988900, 839989800,
    839990700, 839991600, 839992500, 839993400, 839994300, 839995200,
    839996100, 839997000, 839997900, 839998800, 839999700, 840000600,
    840001500, 840002400, 840003300, 840004200, 840005100, 840006000,
    840006900, 840007800, 840008700, 840009600, 840010500, 840011400,
    840012300, 840013200, 840014100, 840015000, 840015900, 840016800,
    840017700, 840018600, 840019500, 840020400, 840021300, 840022200,
    840023100, 840024000, 840024900, 840025800, 840026700, 840027600,
    840028500, 840029400, 840030300, 840031200, 840032100, 840033000,
    840033900, 840034800, 840035700, 840036600, 840037500, 840038400,
    840039300, 840040200, 840041100, 840042000, 840042900, 840043800,
    840044700, 840045600, 840046500, 840047400, 840048300, 840049200,
    840050100, 840051000, 840051900, 840052800, 840053700, 840054600,
    840055500, 840056400, 840057300, 840058200, 840059100, 840060000,
    840060900, 840061800, 840062700, 840063600, 840064500, 840065400,
    840066300, 840067200, 840068100, 840069000, 840069900, 840070800,
    840071700, 840072600, 840073500, 840074400, 840075300, 840076200,
    840077100, 840078000, 840078900, 840079800, 840080700, 840081600,
    840082500, 840083400, 840084300, 840085200, 840086100, 840087000,
    840087900, 840088800, 840089700, 840090600, 840091500, 840092400,
    840093300, 840094200, 840095100, 840096000, 840096900, 840097800,
    840098700, 840099600, 840100500, 840101400, 840102300, 840103200,
    840104100, 840105000, 840105900, 840106800, 840107700, 840108600,
    840109500, 840110400, 840111300, 840112200, 840113100, 840114000,
    840114900, 840115800, 840116700, 840117600, 840118500, 840119400,
    840120300, 840121200, 840122100, 840123000, 840123900, 840124800,
    840125700, 840126600, 840127500, 840128400, 840129300, 840130200,
    840131100, 840132000, 840132900, 840133800, 840134700, 840135600,
    840136500, 840137400, 840138300, 840139200, 840140100, 840141000,
    840141900, 840142800, 840143700, 840144600, 840145500, 840146400,
    840147300, 840148200, 840149100, 840150000, 840150900, 840151800,
    840152700, 840153600, 840154500, 840155400, 840156300, 840157200,
    840158100, 840159000, 840159900, 840160800, 840161700, 840162600,
    840163500, 840164400, 840165300, 840166200, 840167100, 840168000,
    840168900, 840169800, 840170700, 840171600, 840172500, 840173400,
    840174300, 840175200, 840176100, 840177000, 840177900, 840178800,
    840179700, 840180600, 840181500, 840182400, 840183300, 840184200,
    840185100, 840186000, 840186900, 840187800, 840188700, 840189600,
    840190500, 840191400, 840192300, 840193200, 840194100, 840195000,
    840195900, 840196800, 840197700, 840198600, 840199500, 840200400,
    840201300, 840202200, 840203100, 840204000, 840204900, 840205800,
    840206700, 840207600, 840208500, 840209400, 840210300, 840211200,
    840212100, 840213000, 840213900, 840214800, 840215700, 840216600,
    840217500, 840218400, 840219300, 840220200, 840221100, 840222000,
    840222900, 840223800, 840224700, 840225600, 840226500, 840227400,
    840228300, 840229200, 840230100, 840231000, 840231900, 840232800,
    840233700, 840234600, 840235500, 840236400, 840237300, 840238200,
    840239100, 840240000, 840240900, 840241800, 840242700, 840243600,
    840244500, 840245400, 840246300, 840247200, 840248100, 840249000,
    840249900, 840250800, 840251700, 840252600, 840253500, 840254400,
    840255300, 840256200, 840257100, 840258000, 840258900, 840259800,
    840260700, 840261600, 840262500, 840263400, 840264300, 840265200,
    840266100, 840267000, 840267900, 840268800, 840269700, 840270600,
    840271500, 840272400, 840273300, 840274200, 840275100, 840276000,
    840276900, 840277800, 840278700, 840279600, 840280500, 840281400,
    840282300, 840283200, 840284100, 840285000, 840285900, 840286800,
    840287700, 840288600, 840289500, 840290400, 840291300, 840292200,
    840293100, 840294000, 840294900, 840295800, 840296700, 840297600,
    840298500, 840299400, 840300300, 840301200, 840302100, 840303000,
    840303900, 840304800, 840305700, 840306600, 840307500, 840308400,
    840309300, 840310200, 840311100, 840312000, 840312900, 840313800,
    840314700, 840315600, 840316500, 840317400, 840318300, 840319200,
    840320100, 840321000, 840321900, 840322800, 840323700, 840324600,
    840325500, 840326400, 840327300, 840328200, 840329100, 840330000,
    840330900, 840331800, 840332700, 840333600, 840334500, 840335400,
    840336300, 840337200, 840338100, 840339000, 840339900, 840340800,
    840341700, 840342600, 840343500, 840344400, 840345300, 840346200,
    840347100, 840348000, 840348900, 840349800, 840350700, 840351600,
    840352500, 840353400, 840354300, 840355200, 840356100, 840357000,
    840357900, 840358800, 840359700, 840360600, 840361500, 840362400,
    840363300, 840364200, 840365100, 840366000, 840366900, 840367800,
    840368700, 840369600, 840370500, 840371400, 840372300, 840373200,
    840374100, 840375000, 840375900, 840376800, 840377700, 840378600,
    840379500, 840380400, 840381300, 840382200, 840383100, 840384000,
    840384900, 840385800, 840386700, 840387600, 840388500, 840389400,
    840390300, 840391200, 840392100, 840393000, 840393900, 840394800,
    840395700, 840396600, 840397500, 840398400, 840399300, 840400200,
    840401100, 840402000, 840402900, 840403800, 840404700, 840405600,
    840406500, 840407400, 840408300, 840409200, 840410100, 840411000,
    840411900, 840412800, 840413700, 840414600, 840415500, 840416400,
    840417300, 840418200, 840419100, 840420000, 840420900, 840421800,
    840422700, 840423600, 840424500, 840425400, 840426300, 840427200,
    840428100, 840429000, 840429900, 840430800, 840431700, 840432600,
    840433500, 840434400, 840435300, 840436200, 840437100, 840438000,
    840438900, 840439800, 840440700, 840441600, 840442500, 840443400,
    840444300, 840445200, 840446100, 840447000, 840447900, 840448800,
    840449700, 840450600, 840451500, 840452400, 840453300, 840454200,
    840455100, 840456000, 840456900, 840457800, 840458700, 840459600,
    840460500, 840461400, 840462300, 840463200, 840464100, 840465000,
    840465900, 840466800, 840467700, 840468600, 840469500, 840470400,
    840471300, 840472200, 840473100, 840474000, 840474900, 840475800,
    840476700, 840477600, 840478500, 840479400, 840480300, 840481200,
    840482100, 840483000, 840483900, 840484800, 840485700, 840486600,
    840487500, 840488400, 840489300, 840490200, 840491100, 840492000,
    840492900, 840493800, 840494700, 840495600, 840496500, 840497400,
    840498300, 840499200, 840500100, 840501000, 840501900, 840502800,
    840503700, 840504600, 840505500, 840506400, 840507300, 840508200,
    840509100, 840510000, 840510900, 840511800, 840512700, 840513600,
    840514500, 840515400, 840516300, 840517200, 840518100, 840519000,
    840519900, 840520800, 840521700, 840522600, 840523500, 840524400,
    840525300, 840526200, 840527100, 840528000, 840528900, 840529800,
    840530700, 840531600, 840532500, 840533400, 840534300, 840535200,
    840536100, 840537000, 840537900, 840538800, 840539700, 840540600,
    840541500, 840542400, 840543300, 840544200, 840545100, 840546000,
    840546900, 840547800, 840548700, 840549600, 840550500, 840551400,
    840552300, 840553200, 840554100, 840555000, 840555900, 840556800,
    840557700, 840558600, 840559500, 840560400, 840561300, 840562200,
    840563100, 840564000, 840564900, 840565800, 840566700, 840567600,
    840568500, 840569400, 840570300, 840571200, 840572100, 840573000,
    840573900, 840574800, 840575700, 840576600, 840577500, 840578400,
    840579300, 840580200, 840581100, 840582000, 840582900, 840583800,
    840584700, 840585600, 840586500, 840587400, 840588300, 840589200,
    840590100, 840591000, 840591900, 840592800, 840593700, 840594600,
    840595500, 840596400, 840597300, 840598200, 840599100, 840600000,
    840600900, 840601800, 840602700, 840603600, 840604500, 840605400,
    840606300, 840607200, 840608100, 840609000, 840609900, 840610800,
    840611700, 840612600, 840613500, 840614400, 840615300, 840616200,
    840617100, 840618000, 840618900, 840619800, 840620700, 840621600,
    840622500, 840623400, 840624300, 840625200, 840626100, 840627000,
    840627900, 840628800, 840629700, 840630600, 840631500, 840632400,
    840633300, 840634200, 840635100, 840636000, 840636900, 840637800,
    840638700, 840639600, 840640500, 840641400, 840642300, 840643200,
    840644100, 840645000, 840645900, 840646800, 840647700, 840648600,
    840649500, 840650400, 840651300, 840652200, 840653100, 840654000,
    840654900, 840655800, 840656700, 840657600, 840658500, 840659400,
    840660300, 840661200, 840662100, 840663000, 840663900, 840664800,
    840665700, 840666600, 840667500, 840668400, 840669300, 840670200,
    840671100, 840672000, 840672900, 840673800, 840674700, 840675600,
    840676500, 840677400, 840678300, 840679200, 840680100, 840681000,
    840681900, 840682800, 840683700, 840684600, 840685500, 840686400,
    840687300, 840688200, 840689100, 840690000, 840690900, 840691800,
    840692700, 840693600, 840694500, 840695400, 840696300, 840697200,
    840698100, 840699000, 840699900, 840700800, 840701700, 840702600,
    840703500, 840704400, 840705300, 840706200, 840707100, 840708000,
    840708900, 840709800, 840710700, 840711600, 840712500, 840713400,
    840714300, 840715200, 840716100, 840717000, 840717900, 840718800,
    840719700, 840720600, 840721500, 840722400, 840723300, 840724200,
    840725100, 840726000, 840726900, 840727800, 840728700, 840729600,
    840730500, 840731400, 840732300, 840733200, 840734100, 840735000,
    840735900, 840736800, 840737700, 840738600, 840739500, 840740400,
    840741300, 840742200, 840743100, 840744000, 840744900, 840745800,
    840746700, 840747600, 840748500, 840749400, 840750300, 840751200,
    840752100, 840753000, 840753900, 840754800, 840755700, 840756600,
    840757500, 840758400, 840759300, 840760200, 840761100, 840762000,
    840762900, 840763800, 840764700, 840765600, 840766500, 840767400,
    840768300, 840769200, 840770100, 840771000, 840771900, 840772800,
    840773700, 840774600, 840775500, 840776400, 840777300, 840778200,
    840779100, 840780000, 840780900, 840781800, 840782700, 840783600,
    840784500, 840785400, 840786300, 840787200, 840788100, 840789000,
    840789900, 840790800, 840791700, 840792600, 840793500, 840794400,
    840795300, 840796200, 840797100, 840798000, 840798900, 840799800,
    840800700, 840801600, 840802500, 840803400, 840804300, 840805200,
    840806100, 840807000, 840807900, 840808800, 840809700, 840810600,
    840811500, 840812400, 840813300, 840814200, 840815100, 840816000,
    840816900, 840817800, 840818700, 840819600, 840820500, 840821400,
    840822300, 840823200, 840824100, 840825000, 840825900, 840826800,
    840827700, 840828600, 840829500, 840830400, 840831300, 840832200,
    840833100, 840834000, 840834900, 840835800, 840836700, 840837600,
    840838500, 840839400, 840840300, 840841200, 840842100, 840843000,
    840843900, 840844800, 840845700, 840846600, 840847500, 840848400,
    840849300, 840850200, 840851100, 840852000, 840852900, 840853800,
    840854700, 840855600, 840856500, 840857400, 840858300, 840859200,
    840860100, 840861000, 840861900, 840862800, 840863700, 840864600,
    840865500, 840866400, 840867300, 840868200, 840869100, 840870000,
    840870900, 840871800, 840872700, 840873600, 840874500, 840875400,
    840876300, 840877200, 840878100, 840879000, 840879900, 840880800,
    840881700, 840882600, 840883500, 840884400, 840885300, 840886200,
    840887100, 840888000, 840888900, 840889800, 840890700, 840891600,
    840892500, 840893400, 840894300, 840895200, 840896100, 840897000,
    840897900, 840898800, 840899700, 840900600, 840901500, 840902400,
    840903300, 840904200, 840905100, 840906000, 840906900, 840907800,
    840908700, 840909600, 840910500, 840911400, 840912300, 840913200,
    840914100, 840915000, 840915900, 840916800, 840917700, 840918600,
    840919500, 840920400, 840921300, 840922200, 840923100, 840924000,
    840924900, 840925800, 840926700, 840927600, 840928500, 840929400,
    840930300, 840931200, 840932100, 840933000, 840933900, 840934800,
    840935700, 840936600, 840937500, 840938400, 840939300, 840940200,
    840941100, 840942000, 840942900, 840943800, 840944700, 840945600,
    840946500, 840947400, 840948300, 840949200, 840950100, 840951000,
    840951900, 840952800, 840953700, 840954600, 840955500, 840956400,
    840957300, 840958200, 840959100, 840960000, 840960900, 840961800,
    840962700, 840963600, 840964500, 840965400, 840966300, 840967200,
    840968100, 840969000, 840969900, 840970800, 840971700, 840972600,
    840973500, 840974400, 840975300, 840976200, 840977100, 840978000,
    840978900, 840979800, 840980700, 840981600, 840982500, 840983400,
    840984300, 840985200, 840986100, 840987000, 840987900, 840988800,
    840989700, 840990600, 840991500, 840992400, 840993300, 840994200,
    840995100, 840996000, 840996900, 840997800, 840998700, 840999600,
    841000500, 841001400, 841002300, 841003200, 841004100, 841005000,
    841005900, 841006800, 841007700, 841008600, 841009500, 841010400,
    841011300, 841012200, 841013100, 841014000, 841014900, 841015800,
    841016700, 841017600, 841018500, 841019400, 841020300, 841021200,
    841022100, 841023000, 841023900, 841024800, 841025700, 841026600,
    841027500, 841028400, 841029300, 841030200, 841031100, 841032000,
    841032900, 841033800, 841034700, 841035600, 841036500, 841037400,
    841038300, 841039200, 841040100, 841041000, 841041900, 841042800,
    841043700, 841044600, 841045500, 841046400, 841047300, 841048200,
    841049100, 841050000, 841050900, 841051800, 841052700, 841053600,
    841054500, 841055400, 841056300, 841057200, 841058100, 841059000,
    841059900, 841060800, 841061700, 841062600, 841063500, 841064400,
    841065300, 841066200, 841067100, 841068000, 841068900, 841069800,
    841070700, 841071600, 841072500, 841073400, 841074300, 841075200,
    841076100, 841077000, 841077900, 841078800, 841079700, 841080600,
    841081500, 841082400, 841083300, 841084200, 841085100, 841086000,
    841086900, 841087800, 841088700, 841089600, 841090500, 841091400,
    841092300, 841093200, 841094100, 841095000, 841095900, 841096800,
    841097700, 841098600, 841099500, 841100400, 841101300, 841102200,
    841103100, 841104000, 841104900, 841105800, 841106700, 841107600,
    841108500, 841109400, 841110300, 841111200, 841112100, 841113000,
    841113900, 841114800, 841115700, 841116600, 841117500, 841118400,
    841119300, 841120200, 841121100, 841122000, 841122900, 841123800,
    841124700, 841125600, 841126500, 841127400, 841128300, 841129200,
    841130100, 841131000, 841131900, 841132800, 841133700, 841134600,
    841135500, 841136400, 841137300, 841138200, 841139100, 841140000,
    841140900, 841141800, 841142700, 841143600, 841144500, 841145400,
    841146300, 841147200, 841148100, 841149000, 841149900, 841150800,
    841151700, 841152600, 841153500, 841154400, 841155300, 841156200,
    841157100, 841158000, 841158900, 841159800, 841160700, 841161600,
    841162500, 841163400, 841164300, 841165200, 841166100, 841167000,
    841167900, 841168800, 841169700, 841170600, 841171500, 841172400,
    841173300, 841174200, 841175100, 841176000, 841176900, 841177800,
    841178700, 841179600, 841180500, 841181400, 841182300, 841183200,
    841184100, 841185000, 841185900, 841186800, 841187700, 841188600,
    841189500, 841190400, 841191300, 841192200, 841193100, 841194000,
    841194900, 841195800, 841196700, 841197600, 841198500, 841199400,
    841200300, 841201200, 841202100, 841203000, 841203900, 841204800,
    841205700, 841206600, 841207500, 841208400, 841209300, 841210200,
    841211100, 841212000, 841212900, 841213800, 841214700, 841215600,
    841216500, 841217400, 841218300, 841219200, 841220100, 841221000,
    841221900, 841222800, 841223700, 841224600, 841225500, 841226400,
    841227300, 841228200, 841229100, 841230000, 841230900, 841231800,
    841232700, 841233600, 841234500, 841235400, 841236300, 841237200,
    841238100, 841239000, 841239900, 841240800, 841241700, 841242600,
    841243500, 841244400, 841245300, 841246200, 841247100, 841248000,
    841248900, 841249800, 841250700, 841251600, 841252500, 841253400,
    841254300, 841255200, 841256100, 841257000, 841257900, 841258800,
    841259700, 841260600, 841261500, 841262400, 841263300, 841264200,
    841265100, 841266000, 841266900, 841267800, 841268700, 841269600,
    841270500, 841271400, 841272300, 841273200, 841274100, 841275000,
    841275900, 841276800, 841277700, 841278600, 841279500, 841280400,
    841281300, 841282200, 841283100, 841284000, 841284900, 841285800,
    841286700, 841287600, 841288500, 841289400, 841290300, 841291200,
    841292100, 841293000, 841293900, 841294800, 841295700, 841296600,
    841297500, 841298400, 841299300, 841300200, 841301100, 841302000,
    841302900, 841303800, 841304700, 841305600, 841306500, 841307400,
    841308300, 841309200, 841310100, 841311000, 841311900, 841312800,
    841313700, 841314600, 841315500, 841316400, 841317300, 841318200,
    841319100, 841320000, 841320900, 841321800, 841322700, 841323600,
    841324500, 841325400, 841326300, 841327200, 841328100, 841329000,
    841329900, 841330800, 841331700, 841332600, 841333500, 841334400,
    841335300, 841336200, 841337100, 841338000, 841338900, 841339800,
    841340700, 841341600, 841342500, 841343400, 841344300, 841345200,
    841346100, 841347000, 841347900, 841348800, 841349700, 841350600,
    841351500, 841352400, 841353300, 841354200, 841355100, 841356000,
    841356900, 841357800, 841358700, 841359600, 841360500, 841361400,
    841362300, 841363200, 841364100, 841365000, 841365900, 841366800,
    841367700, 841368600, 841369500, 841370400, 841371300, 841372200,
    841373100, 841374000, 841374900, 841375800, 841376700, 841377600,
    841378500, 841379400, 841380300, 841381200, 841382100, 841383000,
    841383900, 841384800, 841385700, 841386600, 841387500, 841388400,
    841389300, 841390200, 841391100, 841392000, 841392900, 841393800,
    841394700, 841395600, 841396500, 841397400, 841398300, 841399200,
    841400100, 841401000, 841401900, 841402800, 841403700, 841404600,
    841405500, 841406400, 841407300, 841408200, 841409100, 841410000,
    841410900, 841411800, 841412700, 841413600, 841414500, 841415400,
    841416300, 841417200, 841418100, 841419000, 841419900, 841420800,
    841421700, 841422600, 841423500, 841424400, 841425300, 841426200,
    841427100, 841428000, 841428900, 841429800, 841430700, 841431600,
    841432500, 841433400, 841434300, 841435200, 841436100, 841437000,
    841437900, 841438800, 841439700, 841440600, 841441500, 841442400,
    841443300, 841444200, 841445100, 841446000, 841446900, 841447800,
    841448700, 841449600, 841450500, 841451400, 841452300, 841453200,
    841454100, 841455000, 841455900, 841456800, 841457700, 841458600,
    841459500, 841460400, 841461300, 841462200, 841463100, 841464000,
    841464900, 841465800, 841466700, 841467600, 841468500, 841469400,
    841470300, 841471200, 841472100, 841473000, 841473900, 841474800,
    841475700, 841476600, 841477500, 841478400, 841479300, 841480200,
    841481100, 841482000, 841482900, 841483800, 841484700, 841485600,
    841486500, 841487400, 841488300, 841489200, 841490100, 841491000,
    841491900, 841492800, 841493700, 841494600, 841495500, 841496400,
    841497300, 841498200, 841499100, 841500000, 841500900, 841501800,
    841502700, 841503600, 841504500, 841505400, 841506300, 841507200,
    841508100, 841509000, 841509900, 841510800, 841511700, 841512600,
    841513500, 841514400, 841515300, 841516200, 841517100, 841518000,
    841518900, 841519800, 841520700, 841521600, 841522500, 841523400,
    841524300, 841525200, 841526100, 841527000, 841527900, 841528800,
    841529700, 841530600, 841531500, 841532400, 841533300, 841534200,
    841535100, 841536000, 841536900, 841537800, 841538700, 841539600,
    841540500, 841541400, 841542300, 841543200, 841544100, 841545000,
    841545900, 841546800, 841547700, 841548600, 841549500, 841550400,
    841551300, 841552200, 841553100, 841554000, 841554900, 841555800,
    841556700, 841557600, 841558500, 841559400, 841560300, 841561200,
    841562100, 841563000, 841563900, 841564800, 841565700, 841566600,
    841567500, 841568400, 841569300, 841570200, 841571100, 841572000,
    841572900, 841573800, 841574700, 841575600, 841576500, 841577400,
    841578300, 841579200, 841580100, 841581000, 841581900, 841582800,
    841583700, 841584600, 841585500, 841586400, 841587300, 841588200,
    841589100, 841590000, 841590900, 841591800, 841592700, 841593600,
    841594500, 841595400, 841596300, 841597200, 841598100, 841599000,
    841599900, 841600800, 841601700, 841602600, 841603500, 841604400,
    841605300, 841606200, 841607100, 841608000, 841608900, 841609800,
    841610700, 841611600, 841612500, 841613400, 841614300, 841615200,
    841616100, 841617000, 841617900, 841618800, 841619700, 841620600,
    841621500, 841622400, 841623300, 841624200, 841625100, 841626000,
    841626900, 841627800, 841628700, 841629600, 841630500, 841631400,
    841632300, 841633200, 841634100, 841635000, 841635900, 841636800,
    841637700, 841638600, 841639500, 841640400, 841641300, 841642200,
    841643100, 841644000, 841644900, 841645800, 841646700, 841647600,
    841648500, 841649400, 841650300, 841651200, 841652100, 841653000,
    841653900, 841654800, 841655700, 841656600, 841657500, 841658400,
    841659300, 841660200, 841661100, 841662000, 841662900, 841663800,
    841664700, 841665600, 841666500, 841667400, 841668300, 841669200,
    841670100, 841671000, 841671900, 841672800, 841673700, 841674600,
    841675500, 841676400, 841677300, 841678200, 841679100, 841680000,
    841680900, 841681800, 841682700, 841683600, 841684500, 841685400,
    841686300, 841687200, 841688100, 841689000, 841689900, 841690800,
    841691700, 841692600, 841693500, 841694400, 841695300, 841696200,
    841697100, 841698000, 841698900, 841699800, 841700700, 841701600,
    841702500, 841703400, 841704300, 841705200, 841706100, 841707000,
    841707900, 841708800, 841709700, 841710600, 841711500, 841712400,
    841713300, 841714200, 841715100, 841716000, 841716900, 841717800,
    841718700, 841719600, 841720500, 841721400, 841722300, 841723200,
    841724100, 841725000, 841725900, 841726800, 841727700, 841728600,
    841729500, 841730400, 841731300, 841732200, 841733100, 841734000,
    841734900, 841735800, 841736700, 841737600, 841738500, 841739400,
    841740300, 841741200, 841742100, 841743000, 841743900, 841744800,
    841745700, 841746600, 841747500, 841748400, 841749300, 841750200,
    841751100, 841752000, 841752900, 841753800, 841754700, 841755600,
    841756500, 841757400, 841758300, 841759200, 841760100, 841761000,
    841761900, 841762800, 841763700, 841764600, 841765500, 841766400,
    841767300, 841768200, 841769100, 841770000, 841770900, 841771800,
    841772700, 841773600, 841774500, 841775400, 841776300, 841777200,
    841778100, 841779000, 841779900, 841780800, 841781700, 841782600,
    841783500, 841784400, 841785300, 841786200, 841787100, 841788000,
    841788900, 841789800, 841790700, 841791600, 841792500, 841793400,
    841794300, 841795200, 841796100, 841797000, 841797900, 841798800,
    841799700, 841800600, 841801500, 841802400, 841803300, 841804200,
    841805100, 841806000, 841806900, 841807800, 841808700, 841809600,
    841810500, 841811400, 841812300, 841813200, 841814100, 841815000,
    841815900, 841816800, 841817700, 841818600, 841819500, 841820400,
    841821300, 841822200, 841823100, 841824000, 841824900, 841825800,
    841826700, 841827600, 841828500, 841829400, 841830300, 841831200,
    841832100, 841833000, 841833900, 841834800, 841835700, 841836600,
    841837500, 841838400, 841839300, 841840200, 841841100, 841842000,
    841842900, 841843800, 841844700, 841845600, 841846500, 841847400,
    841848300, 841849200, 841850100, 841851000, 841851900, 841852800,
    841853700, 841854600, 841855500, 841856400, 841857300, 841858200,
    841859100, 841860000, 841860900, 841861800, 841862700, 841863600,
    841864500, 841865400, 841866300, 841867200, 841868100, 841869000,
    841869900, 841870800, 841871700, 841872600, 841873500, 841874400,
    841875300, 841876200, 841877100, 841878000, 841878900, 841879800,
    841880700, 841881600, 841882500, 841883400, 841884300, 841885200,
    841886100, 841887000, 841887900, 841888800, 841889700, 841890600,
    841891500, 841892400, 841893300, 841894200, 841895100, 841896000,
    841896900, 841897800, 841898700, 841899600, 841900500, 841901400,
    841902300, 841903200, 841904100, 841905000, 841905900, 841906800,
    841907700, 841908600, 841909500, 841910400, 841911300, 841912200,
    841913100, 841914000, 841914900, 841915800, 841916700, 841917600,
    841918500, 841919400, 841920300, 841921200, 841922100, 841923000,
    841923900, 841924800, 841925700, 841926600, 841927500, 841928400,
    841929300, 841930200, 841931100, 841932000, 841932900, 841933800,
    841934700, 841935600, 841936500, 841937400, 841938300, 841939200,
    841940100, 841941000, 841941900, 841942800, 841943700, 841944600,
    841945500, 841946400, 841947300, 841948200, 841949100, 841950000,
    841950900, 841951800, 841952700, 841953600, 841954500, 841955400,
    841956300, 841957200, 841958100, 841959000, 841959900, 841960800,
    841961700, 841962600, 841963500, 841964400, 841965300, 841966200,
    841967100, 841968000, 841968900, 841969800, 841970700, 841971600,
    841972500, 841973400, 841974300, 841975200, 841976100, 841977000,
    841977900, 841978800, 841979700, 841980600, 841981500, 841982400,
    841983300, 841984200, 841985100, 841986000, 841986900, 841987800,
    841988700, 841989600, 841990500, 841991400, 841992300, 841993200,
    841994100, 841995000, 841995900, 841996800, 841997700, 841998600,
    841999500, 842000400, 842001300, 842002200, 842003100, 842004000,
    842004900, 842005800, 842006700, 842007600, 842008500, 842009400,
    842010300, 842011200, 842012100, 842013000, 842013900, 842014800,
    842015700, 842016600, 842017500, 842018400, 842019300, 842020200,
    842021100, 842022000, 842022900, 842023800, 842024700, 842025600,
    842026500, 842027400, 842028300, 842029200, 842030100, 842031000,
    842031900, 842032800, 842033700, 842034600, 842035500, 842036400,
    842037300, 842038200, 842039100, 842040000, 842040900, 842041800,
    842042700, 842043600, 842044500, 842045400, 842046300, 842047200,
    842048100, 842049000, 842049900, 842050800, 842051700, 842052600,
    842053500, 842054400, 842055300, 842056200, 842057100, 842058000,
    842058900, 842059800, 842060700, 842061600, 842062500, 842063400,
    842064300, 842065200, 842066100, 842067000, 842067900, 842068800,
    842069700, 842070600, 842071500, 842072400, 842073300, 842074200,
    842075100, 842076000, 842076900, 842077800, 842078700, 842079600,
    842080500, 842081400, 842082300, 842083200, 842084100, 842085000,
    842085900, 842086800, 842087700, 842088600, 842089500, 842090400,
    842091300, 842092200, 842093100, 842094000, 842094900, 842095800,
    842096700, 842097600, 842098500, 842099400, 842100300, 842101200,
    842102100, 842103000, 842103900, 842104800, 842105700, 842106600,
    842107500, 842108400, 842109300, 842110200, 842111100, 842112000,
    842112900, 842113800, 842114700, 842115600, 842116500, 842117400,
    842118300, 842119200, 842120100, 842121000, 842121900, 842122800,
    842123700, 842124600, 842125500, 842126400, 842127300, 842128200,
    842129100, 842130000, 842130900, 842131800, 842132700, 842133600,
    842134500, 842135400, 842136300, 842137200, 842138100, 842139000,
    842139900, 842140800, 842141700, 842142600, 842143500, 842144400,
    842145300, 842146200, 842147100, 842148000, 842148900, 842149800,
    842150700, 842151600, 842152500, 842153400, 842154300, 842155200,
    842156100, 842157000, 842157900, 842158800, 842159700, 842160600,
    842161500, 842162400, 842163300, 842164200, 842165100, 842166000,
    842166900, 842167800, 842168700, 842169600, 842170500, 842171400,
    842172300, 842173200, 842174100, 842175000, 842175900, 842176800,
    842177700, 842178600, 842179500, 842180400, 842181300, 842182200,
    842183100, 842184000, 842184900, 842185800, 842186700, 842187600,
    842188500, 842189400, 842190300, 842191200, 842192100, 842193000,
    842193900, 842194800, 842195700, 842196600, 842197500, 842198400,
    842199300, 842200200, 842201100, 842202000, 842202900, 842203800,
    842204700, 842205600, 842206500, 842207400, 842208300, 842209200,
    842210100, 842211000, 842211900, 842212800, 842213700, 842214600,
    842215500, 842216400, 842217300, 842218200, 842219100, 842220000,
    842220900, 842221800, 842222700, 842223600, 842224500, 842225400,
    842226300, 842227200, 842228100, 842229000, 842229900, 842230800,
    842231700, 842232600, 842233500, 842234400, 842235300, 842236200,
    842237100, 842238000, 842238900, 842239800, 842240700, 842241600,
    842242500, 842243400, 842244300, 842245200, 842246100, 842247000,
    842247900, 842248800, 842249700, 842250600, 842251500, 842252400,
    842253300, 842254200, 842255100, 842256000, 842256900, 842257800,
    842258700, 842259600, 842260500, 842261400, 842262300, 842263200,
    842264100, 842265000, 842265900, 842266800, 842267700, 842268600,
    842269500, 842270400, 842271300, 842272200, 842273100, 842274000,
    842274900, 842275800, 842276700, 842277600, 842278500, 842279400,
    842280300, 842281200, 842282100, 842283000, 842283900, 842284800,
    842285700, 842286600, 842287500, 842288400, 842289300, 842290200,
    842291100, 842292000, 842292900, 842293800, 842294700, 842295600,
    842296500, 842297400, 842298300, 842299200, 842300100, 842301000,
    842301900, 842302800, 842303700, 842304600, 842305500, 842306400,
    842307300, 842308200, 842309100, 842310000, 842310900, 842311800,
    842312700, 842313600, 842314500, 842315400, 842316300, 842317200,
    842318100, 842319000, 842319900, 842320800, 842321700, 842322600,
    842323500, 842324400, 842325300, 842326200, 842327100, 842328000,
    842328900, 842329800, 842330700, 842331600, 842332500, 842333400,
    842334300, 842335200, 842336100, 842337000, 842337900, 842338800,
    842339700, 842340600, 842341500, 842342400, 842343300, 842344200,
    842345100, 842346000, 842346900, 842347800, 842348700, 842349600,
    842350500, 842351400, 842352300, 842353200, 842354100, 842355000,
    842355900, 842356800, 842357700, 842358600, 842359500, 842360400,
    842361300, 842362200, 842363100, 842364000, 842364900, 842365800,
    842366700, 842367600, 842368500, 842369400, 842370300, 842371200,
    842372100, 842373000, 842373900, 842374800, 842375700, 842376600,
    842377500, 842378400, 842379300, 842380200, 842381100, 842382000,
    842382900, 842383800, 842384700, 842385600, 842386500, 842387400,
    842388300, 842389200, 842390100, 842391000, 842391900, 842392800,
    842393700, 842394600, 842395500, 842396400, 842397300, 842398200,
    842399100, 842400000, 842400900, 842401800, 842402700, 842403600,
    842404500, 842405400, 842406300, 842407200, 842408100, 842409000,
    842409900, 842410800, 842411700, 842412600, 842413500, 842414400,
    842415300, 842416200, 842417100, 842418000, 842418900, 842419800,
    842420700, 842421600, 842422500, 842423400, 842424300, 842425200,
    842426100, 842427000, 842427900, 842428800, 842429700, 842430600,
    842431500, 842432400, 842433300, 842434200, 842435100, 842436000,
    842436900, 842437800, 842438700, 842439600, 842440500, 842441400,
    842442300, 842443200, 842444100, 842445000, 842445900, 842446800,
    842447700, 842448600, 842449500, 842450400, 842451300, 842452200,
    842453100, 842454000, 842454900, 842455800, 842456700, 842457600,
    842458500, 842459400, 842460300, 842461200, 842462100, 842463000,
    842463900, 842464800, 842465700, 842466600, 842467500, 842468400,
    842469300, 842470200, 842471100, 842472000, 842472900, 842473800,
    842474700, 842475600, 842476500, 842477400, 842478300, 842479200,
    842480100, 842481000, 842481900, 842482800, 842483700, 842484600,
    842485500, 842486400, 842487300, 842488200, 842489100, 842490000,
    842490900, 842491800, 842492700, 842493600, 842494500, 842495400,
    842496300, 842497200, 842498100, 842499000, 842499900, 842500800,
    842501700, 842502600, 842503500, 842504400, 842505300, 842506200,
    842507100, 842508000, 842508900, 842509800, 842510700, 842511600,
    842512500, 842513400, 842514300, 842515200, 842516100, 842517000,
    842517900, 842518800, 842519700, 842520600, 842521500, 842522400,
    842523300, 842524200, 842525100, 842526000, 842526900, 842527800,
    842528700, 842529600, 842530500, 842531400, 842532300, 842533200,
    842534100, 842535000, 842535900, 842536800, 842537700, 842538600,
    842539500, 842540400, 842541300, 842542200, 842543100, 842544000,
    842544900, 842545800, 842546700, 842547600, 842548500, 842549400,
    842550300, 842551200, 842552100, 842553000, 842553900, 842554800,
    842555700, 842556600, 842557500, 842558400, 842559300, 842560200,
    842561100, 842562000, 842562900, 842563800, 842564700, 842565600,
    842566500, 842567400, 842568300, 842569200, 842570100, 842571000,
    842571900, 842572800, 842573700, 842574600, 842575500, 842576400,
    842577300, 842578200, 842579100, 842580000, 842580900, 842581800,
    842582700, 842583600, 842584500, 842585400, 842586300, 842587200,
    842588100, 842589000, 842589900, 842590800, 842591700, 842592600,
    842593500, 842594400, 842595300, 842596200, 842597100, 842598000,
    842598900, 842599800, 842600700, 842601600, 842602500, 842603400,
    842604300, 842605200, 842606100, 842607000, 842607900, 842608800,
    842609700, 842610600, 842611500, 842612400, 842613300, 842614200,
    842615100, 842616000, 842616900, 842617800, 842618700, 842619600,
    842620500, 842621400, 842622300, 842623200, 842624100, 842625000,
    842625900, 842626800, 842627700, 842628600, 842629500, 842630400,
    842631300, 842632200, 842633100, 842634000, 842634900, 842635800,
    842636700, 842637600, 842638500, 842639400, 842641200, 842642100,
    842643000, 842643900, 842644800, 842645700, 842646600, 842647500,
    842648400, 842649300, 842650200, 842651100, 842652000, 842652900,
    842653800, 842654700, 842655600, 842656500, 842657400, 842658300,
    842659200, 842660100, 842661000, 842661900, 842662800, 842663700,
    842664600, 842665500, 842666400, 842667300, 842668200, 842669100,
    842670000, 842670900, 842671800, 842672700, 842673600, 842674500,
    842675400, 842676300, 842677200, 842678100, 842679000, 842679900,
    842680800, 842681700, 842682600, 842683500, 842684400, 842685300,
    842686200, 842687100, 842688000, 842688900, 842689800, 842690700,
    842691600, 842692500, 842693400, 842694300, 842695200, 842696100,
    842697000, 842697900, 842698800, 842699700, 842700600, 842701500,
    842702400, 842703300, 842704200, 842705100, 842706000, 842706900,
    842707800, 842708700, 842709600, 842710500, 842711400, 842712300,
    842713200, 842714100, 842715000, 842715900, 842716800, 842717700,
    842718600, 842719500, 842720400, 842721300, 842722200, 842723100,
    842724000, 842724900, 842725800, 842726700, 842727600, 842728500,
    842729400, 842730300, 842731200, 842732100, 842733000, 842733900,
    842734800, 842735700, 842736600, 842737500, 842738400, 842739300,
    842740200, 842741100, 842742000, 842742900, 842743800, 842744700,
    842745600, 842746500, 842747400, 842748300, 842749200, 842750100,
    842751000, 842751900, 842752800, 842753700, 842754600, 842755500,
    842756400, 842757300, 842758200, 842759100, 842760000, 842760900,
    842761800, 842762700, 842763600, 842764500, 842765400, 842766300,
    842767200, 842768100, 842769000, 842769900, 842770800, 842771700,
    842772600, 842773500, 842774400, 842775300, 842776200, 842777100,
    842778000, 842778900, 842779800, 842780700, 842781600, 842782500,
    842783400, 842784300, 842785200, 842786100, 842787000, 842787900,
    842788800, 842789700, 842790600, 842791500, 842792400, 842793300,
    842794200, 842795100, 842796000, 842796900, 842797800, 842798700,
    842799600, 842800500, 842801400, 842802300, 842803200, 842804100,
    842805000, 842805900, 842806800, 842807700, 842808600, 842809500,
    842810400, 842811300, 842812200, 842813100, 842814000, 842814900,
    842815800, 842816700, 842817600, 842818500, 842819400, 842820300,
    842821200, 842822100, 842823000, 842823900, 842824800, 842825700,
    842826600, 842827500, 842828400, 842829300, 842830200, 842831100,
    842832000, 842832900, 842833800, 842834700, 842835600, 842836500,
    842837400, 842838300, 842839200, 842840100, 842841000, 842841900,
    842842800, 842843700, 842844600, 842845500, 842846400, 842847300,
    842848200, 842849100, 842850000, 842850900, 842851800, 842852700,
    842853600, 842854500, 842855400, 842856300, 842857200, 842858100,
    842859000, 842859900, 842860800, 842861700, 842862600, 842863500,
    842864400, 842865300, 842866200, 842867100, 842868000, 842868900,
    842869800, 842870700, 842871600, 842872500, 842873400, 842874300,
    842875200, 842876100, 842877000, 842877900, 842878800, 842879700,
    842880600, 842881500, 842882400, 842883300, 842884200, 842885100,
    842886000, 842886900, 842887800, 842888700, 842889600, 842890500,
    842891400, 842892300, 842893200, 842894100, 842895000, 842895900,
    842896800, 842897700, 842898600, 842899500, 842900400, 842901300,
    842902200, 842903100, 842904000, 842904900, 842905800, 842906700,
    842907600, 842908500, 842909400, 842910300, 842911200, 842912100,
    842913000, 842913900, 842914800, 842915700, 842916600, 842917500,
    842918400, 842919300, 842920200, 842921100, 842922000, 842922900,
    842923800, 842924700, 842925600, 842926500, 842927400, 842928300,
    842929200, 842930100, 842931000, 842931900, 842932800, 842933700,
    842934600, 842935500, 842936400, 842937300, 842938200, 842939100,
    842940000, 842940900, 842941800, 842942700, 842943600, 842944500,
    842945400, 842946300, 842947200, 842948100, 842949000, 842949900,
    842950800, 842951700, 842952600, 842953500, 842954400, 842955300,
    842956200, 842957100, 842958000, 842958900, 842959800, 842960700,
    842961600, 842962500, 842963400, 842964300, 842965200, 842966100,
    842967000, 842967900, 842968800, 842969700, 842970600, 842971500,
    842972400, 842973300, 842974200, 842975100, 842976000, 842976900,
    842977800, 842978700, 842979600, 842980500, 842981400, 842982300,
    842983200, 842984100, 842985000, 842985900, 842986800, 842987700,
    842988600, 842989500, 842990400, 842991300, 842992200, 842993100,
    842994000, 842994900, 842995800, 842996700, 842997600, 842998500,
    842999400, 843000300, 843001200, 843002100, 843003000, 843003900,
    843004800, 843005700, 843006600, 843007500, 843008400, 843009300,
    843010200, 843011100, 843012000, 843012900, 843013800, 843014700,
    843015600, 843016500, 843017400, 843018300, 843019200, 843020100,
    843021000, 843021900, 843022800, 843023700, 843024600, 843025500,
    843026400, 843027300, 843028200, 843029100, 843030000, 843030900,
    843031800, 843032700, 843033600, 843034500, 843035400, 843036300,
    843037200, 843038100, 843039000, 843039900, 843040800, 843041700,
    843042600, 843043500, 843044400, 843045300, 843046200, 843047100,
    843048000, 843048900, 843049800, 843050700, 843051600, 843052500,
    843053400, 843054300, 843055200, 843056100, 843057000, 843057900,
    843058800, 843059700, 843060600, 843061500, 843062400, 843063300,
    843064200, 843065100, 843066000, 843066900, 843067800, 843068700,
    843069600, 843070500, 843071400, 843072300, 843073200, 843074100,
    843075000, 843075900, 843076800, 843077700, 843078600, 843079500,
    843080400, 843081300, 843082200, 843083100, 843084000, 843084900,
    843085800, 843086700, 843087600, 843088500, 843089400, 843090300,
    843091200, 843092100, 843093000, 843093900, 843094800, 843095700,
    843096600, 843097500, 843098400, 843099300, 843100200, 843101100,
    843102000, 843102900, 843103800, 843104700, 843105600, 843106500,
    843107400, 843108300, 843109200, 843110100, 843111000, 843111900,
    843112800, 843113700, 843114600, 843115500, 843116400, 843117300,
    843118200, 843119100, 843120000, 843120900, 843121800, 843122700,
    843123600, 843124500, 843125400, 843126300, 843127200, 843128100,
    843129000, 843129900, 843130800, 843131700, 843132600, 843133500,
    843134400, 843135300, 843136200, 843137100, 843138000, 843138900,
    843139800, 843140700, 843141600, 843142500, 843143400, 843144300,
    843145200, 843146100, 843147000, 843147900, 843148800, 843149700,
    843150600, 843151500, 843152400, 843153300, 843154200, 843155100,
    843156000, 843156900, 843157800, 843158700, 843159600, 843160500,
    843161400, 843162300, 843163200, 843164100, 843165000, 843165900,
    843166800, 843167700, 843168600, 843169500, 843170400, 843171300,
    843172200, 843173100, 843174000, 843174900, 843175800, 843176700,
    843177600, 843178500, 843179400, 843180300, 843181200, 843182100,
    843183000, 843183900, 843184800, 843185700, 843186600, 843187500,
    843188400, 843189300, 843190200, 843191100, 843192000, 843192900,
    843193800, 843194700, 843195600, 843196500, 843197400, 843198300,
    843199200, 843200100, 843201000, 843201900, 843202800, 843203700,
    843204600, 843205500, 843206400, 843207300, 843208200, 843209100,
    843210000, 843210900, 843211800, 843212700, 843213600, 843214500,
    843215400, 843216300, 843217200, 843218100, 843219000, 843219900,
    843220800, 843221700, 843222600, 843223500, 843224400, 843225300,
    843226200, 843227100, 843228000, 843228900, 843229800, 843230700,
    843231600, 843232500, 843233400, 843234300, 843235200, 843236100,
    843237000, 843237900, 843238800, 843239700, 843240600, 843241500,
    843242400, 843243300, 843244200, 843245100, 843246000, 843246900,
    843247800, 843248700, 843249600, 843250500, 843251400, 843252300,
    843253200, 843254100, 843255000, 843255900, 843256800, 843257700,
    843258600, 843259500, 843260400, 843261300, 843262200, 843263100,
    843264000, 843264900, 843265800, 843266700, 843267600, 843268500,
    843269400, 843270300, 843271200, 843272100, 843273000, 843273900,
    843274800, 843275700, 843276600, 843277500, 843278400, 843279300,
    843280200, 843281100, 843282000, 843282900, 843283800, 843284700,
    843285600, 843286500, 843287400, 843288300, 843289200, 843290100,
    843291000, 843291900, 843292800, 843293700, 843294600, 843295500,
    843296400, 843297300, 843298200, 843299100, 843300000, 843300900,
    843301800, 843302700, 843303600, 843304500, 843305400, 843306300,
    843307200, 843308100, 843309000, 843309900, 843310800, 843311700,
    843312600, 843313500, 843314400, 843315300, 843316200, 843317100,
    843318000, 843318900, 843319800, 843320700, 843321600, 843322500,
    843323400, 843324300, 843325200, 843326100, 843327000, 843327900,
    843328800, 843329700, 843330600, 843331500, 843332400, 843333300,
    843334200, 843335100, 843336000, 843336900, 843337800, 843338700,
    843339600, 843340500, 843341400, 843342300, 843343200, 843344100,
    843345000, 843345900, 843346800, 843347700, 843348600, 843349500,
    843350400, 843351300, 843352200, 843353100, 843354000, 843354900,
    843355800, 843356700, 843357600, 843358500, 843359400, 843360300,
    843361200, 843362100, 843363000, 843363900, 843364800, 843365700,
    843366600, 843367500, 843368400, 843369300, 843370200, 843371100,
    843372000, 843372900, 843373800, 843374700, 843375600, 843376500,
    843377400, 843378300, 843379200, 843380100, 843381000, 843381900,
    843382800, 843383700, 843384600, 843385500, 843386400, 843387300,
    843388200, 843389100, 843390000, 843390900, 843391800, 843392700,
    843393600, 843394500, 843395400, 843396300, 843397200, 843398100,
    843399000, 843399900, 843400800, 843401700, 843402600, 843403500,
    843404400, 843405300, 843406200, 843407100, 843408000, 843408900,
    843409800, 843410700, 843411600, 843412500, 843413400, 843414300,
    843415200, 843416100, 843417000, 843417900, 843418800, 843419700,
    843420600, 843421500, 843422400, 843423300, 843424200, 843425100,
    843426000, 843426900, 843427800, 843428700, 843429600, 843430500,
    843431400, 843432300, 843433200, 843434100, 843435000, 843435900,
    843436800, 843437700, 843438600, 843439500, 843440400, 843441300,
    843442200, 843443100, 843444000, 843444900, 843445800, 843446700,
    843447600, 843448500, 843449400, 843450300, 843451200, 843452100,
    843453000, 843453900, 843454800, 843455700, 843456600, 843457500,
    843458400, 843459300, 843460200, 843461100, 843462000, 843462900,
    843463800, 843464700, 843465600, 843466500, 843467400, 843468300,
    843469200, 843470100, 843471000, 843471900, 843472800, 843473700,
    843474600, 843475500, 843476400, 843477300, 843478200, 843479100,
    843480000, 843480900, 843481800, 843482700, 843483600, 843484500,
    843485400, 843486300, 843487200, 843488100, 843489000, 843489900,
    843490800, 843491700, 843492600, 843493500, 843494400, 843495300,
    843496200, 843497100, 843498000, 843498900, 843499800, 843500700,
    843501600, 843502500, 843503400, 843504300, 843505200, 843506100,
    843507000, 843507900, 843508800, 843509700, 843510600, 843511500,
    843512400, 843513300, 843514200, 843515100, 843516000, 843516900,
    843517800, 843518700, 843519600, 843520500, 843521400, 843522300,
    843523200, 843524100, 843525000, 843525900, 843526800, 843527700,
    843528600, 843529500, 843530400, 843531300, 843532200, 843533100,
    843534000, 843534900, 843535800, 843536700, 843537600, 843538500,
    843539400, 843540300, 843541200, 843542100, 843543000, 843543900,
    843544800, 843545700, 843546600, 843547500, 843548400, 843549300,
    843550200, 843551100, 843552000, 843552900, 843553800, 843554700,
    843555600, 843556500, 843557400, 843558300, 843559200, 843560100,
    843561000, 843561900, 843562800, 843563700, 843564600, 843565500,
    843566400, 843567300, 843568200, 843569100, 843570000, 843570900,
    843571800, 843572700, 843573600, 843574500, 843575400, 843576300,
    843577200, 843578100, 843579000, 843579900, 843580800, 843581700,
    843582600, 843583500, 843584400, 843585300, 843586200, 843587100,
    843588000, 843588900, 843589800, 843590700, 843591600, 843592500,
    843593400, 843594300, 843595200, 843596100, 843597000, 843597900,
    843598800, 843599700, 843600600, 843601500, 843602400, 843603300,
    843604200, 843605100, 843606000, 843606900, 843607800, 843608700,
    843609600, 843610500, 843611400, 843612300, 843613200, 843614100,
    843615000, 843615900, 843616800, 843617700, 843618600, 843619500,
    843620400, 843621300, 843622200, 843623100, 843624000, 843624900,
    843625800, 843626700, 843627600, 843628500, 843629400, 843630300,
    843631200, 843632100, 843633000, 843633900, 843634800, 843635700,
    843636600, 843637500, 843638400, 843639300, 843640200, 843641100,
    843642000, 843642900, 843643800, 843644700, 843645600, 843646500,
    843647400, 843648300, 843649200, 843650100, 843651000, 843651900,
    843652800, 843653700, 843654600, 843655500, 843656400, 843657300,
    843658200, 843659100, 843660000, 843660900, 843661800, 843662700,
    843663600, 843664500, 843665400, 843666300, 843667200, 843668100,
    843669000, 843669900, 843670800, 843671700, 843672600, 843673500,
    843674400, 843675300, 843676200, 843677100, 843678000, 843678900,
    843679800, 843680700, 843681600, 843682500, 843683400, 843684300,
    843685200, 843686100, 843687000, 843687900, 843688800, 843689700,
    843690600, 843691500, 843692400, 843693300, 843694200, 843695100,
    843696000, 843696900, 843697800, 843698700, 843699600, 843700500,
    843701400, 843702300, 843703200, 843704100, 843705000, 843705900,
    843706800, 843707700, 843708600, 843709500, 843710400, 843711300,
    843712200, 843713100, 843714000, 843714900, 843715800, 843716700,
    843717600, 843718500, 843719400, 843720300, 843721200, 843722100,
    843723000, 843723900, 843724800, 843725700, 843726600, 843727500,
    843728400, 843729300, 843730200, 843731100, 843732000, 843732900,
    843733800, 843734700, 843735600, 843736500, 843737400, 843738300,
    843739200, 843740100, 843741000, 843741900, 843742800, 843743700,
    843744600, 843745500, 843746400, 843747300, 843748200, 843749100,
    843750000, 843750900, 843751800, 843752700, 843753600, 843754500,
    843755400, 843756300, 843757200, 843758100, 843759000, 843759900,
    843760800, 843761700, 843762600, 843763500, 843764400, 843765300,
    843766200, 843767100, 843768000, 843768900, 843769800, 843770700,
    843771600, 843772500, 843773400, 843774300, 843775200, 843776100,
    843777000, 843777900, 843778800, 843779700, 843780600, 843781500,
    843782400, 843783300, 843784200, 843785100, 843786000, 843786900,
    843787800, 843788700, 843789600, 843790500, 843791400, 843792300,
    843793200, 843794100, 843795000, 843795900, 843796800, 843797700,
    843798600, 843799500, 843800400, 843801300, 843802200, 843803100,
    843804000, 843804900, 843805800, 843806700, 843807600, 843808500,
    843809400, 843810300, 843811200, 843812100, 843813000, 843813900,
    843814800, 843815700, 843816600, 843817500, 843818400, 843819300,
    843820200, 843821100, 843822000, 843822900, 843823800, 843824700,
    843825600, 843826500, 843827400, 843828300, 843829200, 843830100,
    843831000, 843831900, 843832800, 843833700, 843834600, 843835500,
    843836400, 843837300, 843838200, 843839100, 843840000, 843840900,
    843841800, 843842700, 843843600, 843844500, 843845400, 843846300,
    843847200, 843848100, 843849000, 843849900, 843850800, 843851700,
    843852600, 843853500, 843854400, 843855300, 843856200, 843857100,
    843858000, 843858900, 843859800, 843860700, 843861600, 843862500,
    843863400, 843864300, 843865200, 843866100, 843867000, 843867900,
    843868800, 843869700, 843870600, 843871500, 843872400, 843873300,
    843874200, 843875100, 843876000, 843876900, 843877800, 843878700,
    843879600, 843880500, 843881400, 843882300, 843883200, 843884100,
    843885000, 843885900, 843886800, 843887700, 843888600, 843889500,
    843890400, 843891300, 843892200, 843893100, 843894000, 843894900,
    843895800, 843896700, 843897600, 843898500, 843899400, 843900300,
    843901200, 843902100, 843903000, 843903900, 843904800, 843905700,
    843906600, 843907500, 843908400, 843909300, 843910200, 843911100,
    843912000, 843912900, 843913800, 843914700, 843915600, 843916500,
    843917400, 843918300, 843919200, 843920100, 843921000, 843921900,
    843922800, 843923700, 843924600, 843925500, 843926400, 843927300,
    843928200, 843929100, 843930000, 843930900, 843931800, 843932700,
    843933600, 843934500, 843935400, 843936300, 843937200, 843938100,
    843939000, 843939900, 843940800, 843941700, 843942600, 843943500,
    843944400, 843945300, 843946200, 843947100, 843948000, 843948900,
    843949800, 843950700, 843951600, 843952500, 843953400, 843954300,
    843955200, 843956100, 843957000, 843957900, 843958800, 843959700,
    843960600, 843961500, 843962400, 843963300, 843964200, 843965100,
    843966000, 843966900, 843967800, 843968700, 843969600, 843970500,
    843971400, 843972300, 843973200, 843974100, 843975000, 843975900,
    843976800, 843977700, 843978600, 843979500, 843980400, 843981300,
    843982200, 843983100, 843984000, 843984900, 843985800, 843986700,
    843987600, 843988500, 843989400, 843990300, 843991200, 843992100,
    843993000, 843993900, 843994800, 843995700, 843996600, 843997500,
    843998400, 843999300, 844000200, 844001100, 844002000, 844002900,
    844003800, 844004700, 844005600, 844006500, 844007400, 844008300,
    844009200, 844010100, 844011000, 844011900, 844012800, 844013700,
    844014600, 844015500, 844016400, 844017300, 844018200, 844019100,
    844020000, 844020900, 844021800, 844022700, 844023600, 844024500,
    844025400, 844026300, 844027200, 844028100, 844029000, 844029900,
    844030800, 844031700, 844032600, 844033500, 844034400, 844035300,
    844036200, 844037100, 844038000, 844038900, 844039800, 844040700,
    844041600, 844042500, 844043400, 844044300, 844045200, 844046100,
    844047000, 844047900, 844048800, 844049700, 844050600, 844051500,
    844052400, 844053300, 844054200, 844055100, 844056000, 844056900,
    844057800, 844058700, 844059600, 844060500, 844061400, 844062300,
    844063200, 844064100, 844065000, 844065900, 844066800, 844067700,
    844068600, 844069500, 844070400, 844071300, 844072200, 844073100,
    844074000, 844074900, 844075800, 844076700, 844077600, 844078500,
    844079400, 844080300, 844081200, 844082100, 844083000, 844083900,
    844084800, 844085700, 844086600, 844087500, 844088400, 844089300,
    844090200, 844091100, 844092000, 844092900, 844093800, 844094700,
    844095600, 844096500, 844097400, 844098300, 844099200, 844100100,
    844101000, 844101900, 844102800, 844103700, 844104600, 844105500,
    844106400, 844107300, 844108200, 844109100, 844110000, 844110900,
    844111800, 844112700, 844113600, 844114500, 844115400, 844116300,
    844117200, 844118100, 844119000, 844119900, 844120800, 844121700,
    844122600, 844123500, 844124400, 844125300, 844126200, 844127100,
    844128000, 844128900, 844129800, 844130700, 844131600, 844132500,
    844133400, 844134300, 844135200, 844136100, 844137000, 844137900,
    844138800, 844139700, 844140600, 844141500, 844142400, 844143300,
    844144200, 844145100, 844146000, 844146900, 844147800, 844148700,
    844149600, 844150500, 844151400, 844152300, 844153200, 844154100,
    844155000, 844155900, 844156800, 844157700, 844158600, 844159500,
    844160400, 844161300, 844162200, 844163100, 844164000, 844164900,
    844165800, 844166700, 844167600, 844168500, 844169400, 844170300,
    844171200, 844172100, 844173000, 844173900, 844174800, 844175700,
    844176600, 844177500, 844178400, 844179300, 844180200, 844181100,
    844182000, 844182900, 844183800, 844184700, 844185600, 844186500,
    844187400, 844188300, 844189200, 844190100, 844191000, 844191900,
    844192800, 844193700, 844194600, 844195500, 844196400, 844197300,
    844198200, 844199100, 844200000, 844200900, 844201800, 844202700,
    844203600, 844204500, 844205400, 844206300, 844207200, 844208100,
    844209000, 844209900, 844210800, 844211700, 844212600, 844213500,
    844214400, 844215300, 844216200, 844217100, 844218000, 844218900,
    844219800, 844220700, 844221600, 844222500, 844223400, 844224300,
    844225200, 844226100, 844227000, 844227900, 844228800, 844229700,
    844230600, 844231500, 844232400, 844233300, 844234200, 844235100,
    844236000, 844236900, 844237800, 844238700, 844239600, 844240500,
    844241400, 844242300, 844243200, 844244100, 844245000, 844245900,
    844246800, 844247700, 844248600, 844249500, 844250400, 844251300,
    844252200, 844253100, 844254000, 844254900, 844255800, 844256700,
    844257600, 844258500, 844259400, 844260300, 844261200, 844262100,
    844263000, 844263900, 844264800, 844265700, 844266600, 844267500,
    844268400, 844269300, 844270200, 844271100, 844272000, 844272900,
    844273800, 844274700, 844275600, 844276500, 844277400, 844278300,
    844279200, 844280100, 844281000, 844281900, 844282800, 844283700,
    844284600, 844285500, 844286400, 844287300, 844288200, 844289100,
    844290000, 844290900, 844291800, 844292700, 844293600, 844294500,
    844295400, 844296300, 844297200, 844298100, 844299000, 844299900,
    844300800, 844301700, 844302600, 844303500, 844304400, 844305300,
    844306200, 844307100, 844308000, 844308900, 844309800, 844310700,
    844311600, 844312500, 844313400, 844314300, 844315200, 844316100,
    844317000, 844317900, 844318800, 844319700, 844320600, 844321500,
    844322400, 844323300, 844324200, 844325100, 844326000, 844326900,
    844327800, 844328700, 844329600, 844330500, 844331400, 844332300,
    844333200, 844334100, 844335000, 844335900, 844336800, 844337700,
    844338600, 844339500, 844340400, 844341300, 844342200, 844343100,
    844344000, 844344900, 844345800, 844346700, 844347600, 844348500,
    844349400, 844350300, 844351200, 844352100, 844353000, 844353900,
    844354800, 844355700, 844356600, 844357500, 844358400, 844359300,
    844360200, 844361100, 844362000, 844362900, 844363800, 844364700,
    844365600, 844366500, 844367400, 844368300, 844369200, 844370100,
    844371000, 844371900, 844372800, 844373700, 844374600, 844375500,
    844376400, 844377300, 844378200, 844379100, 844380000, 844380900,
    844381800, 844382700, 844383600, 844384500, 844385400, 844386300,
    844387200, 844388100, 844389000, 844389900, 844390800, 844391700,
    844392600, 844393500, 844394400, 844395300, 844396200, 844397100,
    844398000, 844398900, 844399800, 844400700, 844401600, 844402500,
    844403400, 844404300, 844405200, 844406100, 844407000, 844407900,
    844408800, 844409700, 844410600, 844411500, 844412400, 844413300,
    844414200, 844415100, 844416000, 844416900, 844417800, 844418700,
    844419600, 844420500, 844421400, 844422300, 844423200, 844424100,
    844425000, 844425900, 844426800, 844427700, 844428600, 844429500,
    844430400, 844431300, 844432200, 844433100, 844434000, 844434900,
    844435800, 844436700, 844437600, 844438500, 844439400, 844440300,
    844441200, 844442100, 844443000, 844443900, 844444800, 844445700,
    844446600, 844447500, 844448400, 844449300, 844450200, 844451100,
    844452000, 844452900, 844453800, 844454700, 844455600, 844456500,
    844457400, 844458300, 844459200, 844460100, 844461000, 844461900,
    844462800, 844463700, 844464600, 844465500, 844466400, 844467300,
    844468200, 844469100, 844470000, 844470900, 844471800, 844472700,
    844473600, 844474500, 844475400, 844476300, 844477200, 844478100,
    844479000, 844479900, 844480800, 844481700, 844482600, 844483500,
    844484400, 844485300, 844486200, 844487100, 844488000, 844488900,
    844489800, 844490700, 844491600, 844492500, 844493400, 844494300,
    844495200, 844496100, 844497000, 844497900, 844498800, 844499700,
    844500600, 844501500, 844502400, 844503300, 844504200, 844505100,
    844506000, 844506900, 844507800, 844508700, 844509600, 844510500,
    844511400, 844512300, 844513200, 844514100, 844515000, 844515900,
    844516800, 844517700, 844518600, 844519500, 844520400, 844521300,
    844522200, 844523100, 844524000, 844524900, 844525800, 844526700,
    844527600, 844528500, 844529400, 844530300, 844531200, 844532100,
    844533000, 844533900, 844534800, 844535700, 844536600, 844537500,
    844538400, 844539300, 844540200, 844541100, 844542000, 844542900,
    844543800, 844544700, 844545600, 844546500, 844547400, 844548300,
    844549200, 844550100, 844551000, 844551900, 844552800, 844553700,
    844554600, 844555500, 844556400, 844557300, 844558200, 844559100,
    844560000, 844560900, 844561800, 844562700, 844563600, 844564500,
    844565400, 844566300, 844567200, 844568100, 844569000, 844569900,
    844570800, 844571700, 844572600, 844573500, 844574400, 844575300,
    844576200, 844577100, 844578000, 844578900, 844579800, 844580700,
    844581600, 844582500, 844583400, 844584300, 844585200, 844586100,
    844587000, 844587900, 844588800, 844589700, 844590600, 844591500,
    844592400, 844593300, 844594200, 844595100, 844596000, 844596900,
    844597800, 844598700, 844599600, 844600500, 844601400, 844602300,
    844603200, 844604100, 844605000, 844605900, 844606800, 844607700,
    844608600, 844609500, 844610400, 844611300, 844612200, 844613100,
    844614000, 844614900, 844615800, 844616700, 844617600, 844618500,
    844619400, 844620300, 844621200, 844622100, 844623000, 844623900,
    844624800, 844625700, 844626600, 844627500, 844628400, 844629300,
    844630200, 844631100, 844632000, 844632900, 844633800, 844634700,
    844635600, 844636500, 844637400, 844638300, 844639200, 844640100,
    844641000, 844641900, 844642800, 844643700, 844644600, 844645500,
    844646400, 844647300, 844648200, 844649100, 844650000, 844650900,
    844651800, 844652700, 844653600, 844654500, 844655400, 844656300,
    844657200, 844658100, 844659000, 844659900, 844660800, 844661700,
    844662600, 844663500, 844664400, 844665300, 844666200, 844667100,
    844668000, 844668900, 844669800, 844670700, 844671600, 844672500,
    844673400, 844674300, 844675200, 844676100, 844677000, 844677900,
    844678800, 844679700, 844680600, 844681500, 844682400, 844683300,
    844684200, 844685100, 844686000, 844686900, 844687800, 844688700,
    844689600, 844690500, 844691400, 844692300, 844693200, 844694100,
    844695000, 844695900, 844696800, 844697700, 844698600, 844699500,
    844700400, 844701300, 844702200, 844703100, 844704000, 844704900,
    844705800, 844706700, 844707600, 844708500, 844709400, 844710300,
    844711200, 844712100, 844713000, 844713900, 844714800, 844715700,
    844716600, 844717500, 844718400, 844719300, 844720200, 844721100,
    844722000, 844722900, 844723800, 844724700, 844725600, 844726500,
    844727400, 844728300, 844729200, 844731000, 844731900, 844732800,
    844733700, 844734600, 844735500, 844736400, 844737300, 844738200,
    844739100, 844740000, 844740900, 844741800, 844742700, 844743600,
    844744500, 844745400, 844746300, 844747200, 844748100, 844749000,
    844749900, 844750800, 844751700, 844752600, 844753500, 844754400,
    844755300, 844756200, 844757100, 844758000, 844758900, 844759800,
    844760700, 844761600, 844762500, 844763400, 844764300, 844765200,
    844766100, 844767000, 844767900, 844768800, 844769700, 844770600,
    844771500, 844772400, 844773300, 844774200, 844775100, 844776000,
    844776900, 844777800, 844778700, 844779600, 844780500, 844781400,
    844782300, 844783200, 844784100, 844785000, 844785900, 844786800,
    844787700, 844788600, 844789500, 844790400, 844791300, 844792200,
    844793100, 844794000, 844794900, 844795800, 844796700, 844797600,
    844798500, 844799400, 844800300, 844801200, 844802100, 844803000,
    844803900, 844804800, 844805700, 844806600, 844807500, 844808400,
    844809300, 844810200, 844811100, 844812000, 844812900, 844813800,
    844814700, 844815600, 844816500, 844817400, 844818300, 844819200,
    844820100, 844821000, 844821900, 844822800, 844823700, 844824600,
    844825500, 844826400, 844827300, 844828200, 844829100, 844830000,
    844830900, 844831800, 844832700, 844833600, 844834500, 844835400,
    844836300, 844837200, 844838100, 844839000, 844839900, 844840800,
    844841700, 844842600, 844843500, 844844400, 844845300, 844846200,
    844847100, 844848000, 844848900, 844849800, 844850700, 844851600,
    844852500, 844853400, 844854300, 844855200, 844856100, 844857000,
    844857900, 844858800, 844859700, 844860600, 844861500, 844862400,
    844863300, 844864200, 844865100, 844866000, 844866900, 844867800,
    844868700, 844869600, 844870500, 844871400, 844872300, 844873200,
    844874100, 844875000, 844875900, 844876800, 844877700, 844878600,
    844879500, 844880400, 844881300, 844882200, 844883100, 844884000,
    844884900, 844885800, 844886700, 844887600, 844888500, 844889400,
    844890300, 844891200, 844892100, 844893000, 844893900, 844894800,
    844895700, 844896600, 844897500, 844898400, 844899300, 844900200,
    844901100, 844902000, 844902900, 844903800, 844904700, 844905600,
    844906500, 844907400, 844908300, 844909200, 844910100, 844911000,
    844911900, 844912800, 844913700, 844914600, 844915500, 844916400,
    844917300, 844918200, 844919100, 844920000, 844920900, 844921800,
    844922700, 844923600, 844924500, 844925400, 844926300, 844927200,
    844928100, 844929000, 844929900, 844930800, 844931700, 844932600,
    844933500, 844934400, 844935300, 844936200, 844937100, 844938000,
    844938900, 844939800, 844940700, 844941600, 844942500, 844943400,
    844944300, 844945200, 844946100, 844947000, 844947900, 844948800,
    844949700, 844950600, 844951500, 844952400, 844953300, 844954200,
    844955100, 844956000, 844956900, 844957800, 844958700, 844959600,
    844960500, 844961400, 844962300, 844963200, 844964100, 844965000,
    844965900, 844966800, 844967700, 844968600, 844969500, 844970400,
    844971300, 844972200, 844973100, 844974000, 844974900, 844975800,
    844976700, 844977600, 844978500, 844979400, 844980300, 844981200,
    844982100, 844983000, 844983900, 844984800, 844985700, 844986600,
    844987500, 844988400, 844989300, 844990200, 844991100, 844992000,
    844992900, 844993800, 844994700, 844995600, 844996500, 844997400,
    844998300, 844999200, 845000100, 845001000, 845001900, 845002800,
    845003700, 845004600, 845005500, 845006400, 845007300, 845008200,
    845009100, 845010000, 845010900, 845011800, 845012700, 845013600,
    845014500, 845015400, 845016300, 845017200, 845018100, 845019000,
    845019900, 845020800, 845021700, 845022600, 845023500, 845024400,
    845025300, 845026200, 845027100, 845028000, 845028900, 845029800,
    845030700, 845031600, 845032500, 845033400, 845034300, 845035200,
    845036100, 845037000, 845037900, 845038800, 845039700, 845040600,
    845041500, 845042400, 845043300, 845044200, 845045100, 845046000,
    845046900, 845047800, 845048700, 845049600, 845050500, 845051400,
    845052300, 845053200, 845054100, 845055000, 845055900, 845056800,
    845057700, 845058600, 845059500, 845060400, 845061300, 845062200,
    845063100, 845064000, 845064900, 845065800, 845066700, 845067600,
    845068500, 845069400, 845070300, 845071200, 845072100, 845073000,
    845073900, 845074800, 845075700, 845076600, 845077500, 845078400,
    845079300, 845080200, 845081100, 845082000, 845082900, 845083800,
    845084700, 845085600, 845086500, 845087400, 845088300, 845089200,
    845090100, 845091000, 845091900, 845092800, 845093700, 845094600,
    845095500, 845096400, 845097300, 845098200, 845099100, 845100000,
    845100900, 845101800, 845102700, 845103600, 845104500, 845105400,
    845106300, 845107200, 845108100, 845109000, 845109900, 845110800,
    845111700, 845112600, 845113500, 845114400, 845115300, 845116200,
    845117100, 845118000, 845118900, 845119800, 845120700, 845121600,
    845122500, 845123400, 845124300, 845125200, 845126100, 845127000,
    845127900, 845128800, 845129700, 845130600, 845131500, 845132400,
    845133300, 845134200, 845135100, 845136000, 845136900, 845137800,
    845138700, 845139600, 845140500, 845141400, 845142300, 845143200,
    845144100, 845145000, 845145900, 845146800, 845147700, 845148600,
    845149500, 845150400, 845151300, 845152200, 845153100, 845154000,
    845154900, 845155800, 845156700, 845157600, 845158500, 845159400,
    845160300, 845161200, 845162100, 845163000, 845163900, 845164800,
    845165700, 845166600, 845167500, 845168400, 845169300, 845170200,
    845171100, 845172000, 845172900, 845173800, 845174700, 845175600,
    845176500, 845177400, 845178300, 845179200, 845180100, 845181000,
    845181900, 845182800, 845183700, 845184600, 845185500, 845186400,
    845187300, 845188200, 845189100, 845190000, 845190900, 845191800,
    845192700, 845193600, 845194500, 845195400, 845196300, 845197200,
    845198100, 845199000, 845199900, 845200800, 845201700, 845202600,
    845203500, 845204400, 845205300, 845206200, 845207100, 845208000,
    845208900, 845209800, 845210700, 845211600, 845212500, 845213400,
    845214300, 845215200, 845216100, 845217000, 845217900, 845218800,
    845219700, 845220600, 845221500, 845222400, 845223300, 845224200,
    845225100, 845226000, 845226900, 845227800, 845228700, 845229600,
    845230500, 845231400, 845232300, 845233200, 845234100, 845235000,
    845235900, 845236800, 845237700, 845238600, 845239500, 845240400,
    845241300, 845242200, 845243100, 845244000, 845244900, 845245800,
    845246700, 845247600, 845248500, 845249400, 845250300, 845251200,
    845252100, 845253000, 845253900, 845254800, 845255700, 845256600,
    845257500, 845258400, 845259300, 845260200, 845261100, 845262000,
    845262900, 845263800, 845264700, 845265600, 845266500, 845267400,
    845268300, 845269200, 845270100, 845271000, 845271900, 845272800,
    845273700, 845274600, 845275500, 845276400, 845277300, 845278200,
    845279100, 845280000, 845280900, 845281800, 845282700, 845283600,
    845284500, 845285400, 845286300, 845287200, 845288100, 845289000,
    845289900, 845290800, 845291700, 845292600, 845293500, 845294400,
    845295300, 845296200, 845297100, 845298000, 845298900, 845299800,
    845300700, 845301600, 845302500, 845303400, 845304300, 845305200,
    845306100, 845307000, 845307900, 845308800, 845309700, 845310600,
    845311500, 845312400, 845313300, 845314200, 845315100, 845316000,
    845316900, 845317800, 845318700, 845319600, 845320500, 845321400,
    845322300, 845323200, 845324100, 845325000, 845325900, 845326800,
    845327700, 845328600, 845329500, 845330400, 845331300, 845332200,
    845333100, 845334000, 845334900, 845335800, 845336700, 845337600,
    845338500, 845339400, 845340300, 845341200, 845342100, 845343000,
    845343900, 845344800, 845345700, 845346600, 845347500, 845348400,
    845349300, 845350200, 845351100, 845352000, 845352900, 845353800,
    845354700, 845355600, 845356500, 845357400, 845358300, 845359200,
    845360100, 845361000, 845361900, 845362800, 845363700, 845364600,
    845365500, 845366400, 845367300, 845368200, 845369100, 845370000,
    845370900, 845371800, 845372700, 845373600, 845374500, 845375400,
    845376300, 845377200, 845378100, 845379000, 845379900, 845380800,
    845381700, 845382600, 845383500, 845384400, 845385300, 845386200,
    845387100, 845388000, 845388900, 845389800, 845390700, 845391600,
    845392500, 845393400, 845394300, 845395200, 845396100, 845397000,
    845397900, 845398800, 845399700, 845400600, 845401500, 845402400,
    845403300, 845404200, 845405100, 845406000, 845406900, 845407800,
    845408700, 845409600, 845410500, 845411400, 845412300, 845413200,
    845414100, 845415000, 845415900, 845416800, 845417700, 845418600,
    845419500, 845420400, 845421300, 845422200, 845423100, 845424000,
    845424900, 845425800, 845426700, 845427600, 845428500, 845429400,
    845430300, 845431200, 845432100, 845433000, 845433900, 845434800,
    845435700, 845436600, 845437500, 845438400, 845439300, 845440200,
    845441100, 845442000, 845442900, 845443800, 845444700, 845445600,
    845446500, 845447400, 845448300, 845449200, 845450100, 845451000,
    845451900, 845452800, 845453700, 845454600, 845455500, 845456400,
    845457300, 845458200, 845459100, 845460000, 845460900, 845461800,
    845462700, 845463600, 845464500, 845465400, 845466300, 845467200,
    845468100, 845469000, 845469900, 845470800, 845471700, 845472600,
    845473500, 845474400, 845475300, 845476200, 845477100, 845478000,
    845478900, 845479800, 845480700, 845481600, 845482500, 845483400,
    845484300, 845485200, 845486100, 845487000, 845487900, 845488800,
    845489700, 845490600, 845491500, 845492400, 845493300, 845494200,
    845495100, 845496000, 845496900, 845497800, 845498700, 845499600,
    845500500, 845501400, 845502300, 845503200, 845504100, 845505000,
    845505900, 845506800, 845507700, 845508600, 845509500, 845510400,
    845511300, 845512200, 845513100, 845514000, 845514900, 845515800,
    845516700, 845517600, 845518500, 845519400, 845520300, 845521200,
    845522100, 845523000, 845523900, 845524800, 845525700, 845526600,
    845527500, 845528400, 845529300, 845530200, 845531100, 845532000,
    845532900, 845533800, 845534700, 845535600, 845536500, 845537400,
    845538300, 845539200, 845540100, 845541000, 845541900, 845542800,
    845543700, 845544600, 845545500, 845546400, 845547300, 845548200,
    845549100, 845550000, 845550900, 845551800, 845552700, 845553600,
    845554500, 845555400, 845556300, 845557200, 845558100, 845559000,
    845559900, 845560800, 845561700, 845562600, 845563500, 845564400,
    845565300, 845566200, 845567100, 845568000, 845568900, 845569800,
    845570700, 845571600, 845572500, 845573400, 845574300, 845575200,
    845576100, 845577000, 845577900, 845578800, 845579700, 845580600,
    845581500, 845582400, 845583300, 845584200, 845585100, 845586000,
    845586900, 845587800, 845588700, 845589600, 845590500, 845591400,
    845592300, 845593200, 845594100, 845595000, 845595900, 845596800,
    845597700, 845598600, 845599500, 845600400, 845601300, 845602200,
    845603100, 845604000, 845604900, 845605800, 845606700, 845607600,
    845608500, 845609400, 845610300, 845611200, 845612100, 845613000,
    845613900, 845614800, 845615700, 845616600, 845617500, 845618400,
    845619300, 845620200, 845621100, 845622000, 845622900, 845623800,
    845624700, 845625600, 845626500, 845627400, 845628300, 845629200,
    845630100, 845631000, 845631900, 845632800, 845633700, 845634600,
    845635500, 845636400, 845637300, 845638200, 845639100, 845640000,
    845640900, 845641800, 845642700, 845643600, 845644500, 845645400,
    845646300, 845647200, 845648100, 845649000, 845649900, 845650800,
    845651700, 845652600, 845653500, 845654400, 845655300, 845656200,
    845657100, 845658000, 845658900, 845659800, 845660700, 845661600,
    845662500, 845663400, 845664300, 845665200, 845666100, 845667000,
    845667900, 845668800, 845669700, 845670600, 845671500, 845672400,
    845673300, 845674200, 845675100, 845676000, 845676900, 845677800,
    845678700, 845679600, 845680500, 845681400, 845682300, 845683200,
    845684100, 845685000, 845685900, 845686800, 845687700, 845688600,
    845689500, 845690400, 845691300, 845692200, 845693100, 845694000,
    845694900, 845695800, 845696700, 845697600, 845698500, 845699400,
    845700300, 845701200, 845702100, 845703000, 845703900, 845704800,
    845705700, 845706600, 845707500, 845708400, 845709300, 845710200,
    845711100, 845712000, 845712900, 845713800, 845714700, 845715600,
    845716500, 845717400, 845718300, 845719200, 845720100, 845721000,
    845721900, 845722800, 845723700, 845724600, 845725500, 845726400,
    845727300, 845728200, 845729100, 845730000, 845730900, 845731800,
    845732700, 845733600, 845734500, 845735400, 845736300, 845737200,
    845738100, 845739000, 845739900, 845740800, 845741700, 845742600,
    845743500, 845744400, 845745300, 845746200, 845747100, 845748000,
    845748900, 845749800, 845750700, 845751600, 845752500, 845753400,
    845754300, 845755200, 845756100, 845757000, 845757900, 845758800,
    845759700, 845760600, 845761500, 845762400, 845763300, 845764200,
    845765100, 845766000, 845766900, 845767800, 845768700, 845769600,
    845770500, 845771400, 845772300, 845773200, 845774100, 845775000,
    845775900, 845776800, 845777700, 845778600, 845779500, 845780400,
    845781300, 845782200, 845783100, 845784000, 845784900, 845785800,
    845786700, 845787600, 845788500, 845789400, 845790300, 845791200,
    845792100, 845793000, 845793900, 845794800, 845795700, 845796600,
    845797500, 845798400, 845799300, 845800200, 845801100, 845802000,
    845802900, 845803800, 845804700, 845805600, 845806500, 845807400,
    845808300, 845809200, 845810100, 845811000, 845811900, 845812800,
    845813700, 845814600, 845815500, 845816400, 845817300, 845818200,
    845819100, 845820000, 845820900, 845821800, 845822700, 845823600,
    845824500, 845825400, 845826300, 845827200, 845828100, 845829000,
    845829900, 845830800, 845831700, 845832600, 845833500, 845834400,
    845835300, 845836200, 845837100, 845838000, 845838900, 845839800,
    845840700, 845841600, 845842500, 845843400, 845844300, 845845200,
    845846100, 845847000, 845847900, 845848800, 845849700, 845850600,
    845851500, 845852400, 845853300, 845854200, 845855100, 845856000,
    845856900, 845857800, 845858700, 845859600, 845860500, 845861400,
    845862300, 845863200, 845864100, 845865000, 845865900, 845866800,
    845867700, 845868600, 845869500, 845870400, 845871300, 845872200,
    845873100, 845874000, 845874900, 845875800, 845876700, 845877600,
    845878500, 845879400, 845880300, 845881200, 845882100, 845883000,
    845883900, 845884800, 845885700, 845886600, 845887500, 845888400,
    845889300, 845890200, 845891100, 845892000, 845892900, 845893800,
    845894700, 845895600, 845896500, 845897400, 845898300, 845899200,
    845900100, 845901000, 845901900, 845902800, 845903700, 845904600,
    845905500, 845906400, 845907300, 845908200, 845909100, 845910000,
    845910900, 845911800, 845912700, 845913600, 845914500, 845915400,
    845916300, 845917200, 845918100, 845919000, 845919900, 845920800,
    845921700, 845922600, 845923500, 845924400, 845925300, 845926200,
    845927100, 845928000, 845928900, 845929800, 845930700, 845931600,
    845932500, 845933400, 845934300, 845935200, 845936100, 845937000,
    845937900, 845938800, 845939700, 845940600, 845941500, 845942400,
    845943300, 845944200, 845945100, 845946000, 845946900, 845947800,
    845948700, 845949600, 845950500, 845951400, 845952300, 845953200,
    845954100, 845955000, 845955900, 845956800, 845957700, 845958600,
    845959500, 845960400, 845961300, 845962200, 845963100, 845964000,
    845964900, 845965800, 845966700, 845967600, 845968500, 845969400,
    845970300, 845971200, 845972100, 845973000, 845973900, 845974800,
    845975700, 845976600, 845977500, 845978400, 845979300, 845980200,
    845981100, 845982000, 845982900, 845983800, 845984700, 845985600,
    845986500, 845987400, 845988300, 845989200, 845990100, 845991000,
    845991900, 845992800, 845993700, 845994600, 845995500, 845996400,
    845997300, 845998200, 845999100, 846000000, 846000900, 846001800,
    846002700, 846003600, 846004500, 846005400, 846006300, 846007200,
    846008100, 846009000, 846009900, 846010800, 846011700, 846012600,
    846013500, 846014400, 846015300, 846016200, 846017100, 846018000,
    846018900, 846019800, 846020700, 846021600, 846022500, 846023400,
    846024300, 846025200, 846026100, 846027000, 846027900, 846028800,
    846029700, 846030600, 846031500, 846032400, 846033300, 846034200,
    846035100, 846036000, 846036900, 846037800, 846038700, 846039600,
    846040500, 846041400, 846042300, 846043200, 846044100, 846045000,
    846045900, 846046800, 846047700, 846048600, 846049500, 846050400,
    846051300, 846052200, 846053100, 846054000, 846054900, 846055800,
    846056700, 846057600, 846058500, 846059400, 846060300, 846061200,
    846062100, 846063000, 846063900, 846064800, 846065700, 846066600,
    846067500, 846068400, 846069300, 846070200, 846071100, 846072000,
    846072900, 846073800, 846074700, 846075600, 846076500, 846077400,
    846078300, 846079200, 846080100, 846081000, 846081900, 846082800,
    846083700, 846084600, 846085500, 846086400, 846087300, 846088200,
    846089100, 846090000, 846090900, 846091800, 846092700, 846093600,
    846094500, 846095400, 846096300, 846097200, 846098100, 846099000,
    846099900, 846100800, 846101700, 846102600, 846103500, 846104400,
    846105300, 846106200, 846107100, 846108000, 846108900, 846109800,
    846110700, 846111600, 846112500, 846113400, 846114300, 846115200,
    846116100, 846117000, 846117900, 846118800, 846119700, 846120600,
    846121500, 846122400, 846123300, 846124200, 846125100, 846126000,
    846126900, 846127800, 846128700, 846129600, 846130500, 846131400,
    846132300, 846133200, 846134100, 846135000, 846135900, 846136800,
    846137700, 846138600, 846139500, 846140400, 846141300, 846142200,
    846143100, 846144000, 846144900, 846145800, 846146700, 846147600,
    846148500, 846149400, 846150300, 846151200, 846152100, 846153000,
    846153900, 846154800, 846155700, 846156600, 846157500, 846158400,
    846159300, 846160200, 846161100, 846162000, 846162900, 846163800,
    846164700, 846165600, 846166500, 846167400, 846168300, 846169200,
    846170100, 846171000, 846171900, 846172800, 846173700, 846174600,
    846175500, 846176400, 846177300, 846178200, 846179100, 846180000,
    846180900, 846181800, 846182700, 846183600, 846184500, 846185400,
    846186300, 846187200, 846188100, 846189000, 846189900, 846190800,
    846191700, 846192600, 846193500, 846194400, 846195300, 846196200,
    846197100, 846198000, 846198900, 846199800, 846200700, 846201600,
    846202500, 846203400, 846204300, 846205200, 846206100, 846207000,
    846207900, 846208800, 846209700, 846210600, 846211500, 846212400,
    846213300, 846214200, 846215100, 846216000, 846216900, 846217800,
    846218700, 846219600, 846220500, 846221400, 846222300, 846223200,
    846224100, 846225000, 846225900, 846226800, 846227700, 846228600,
    846229500, 846230400, 846231300, 846232200, 846233100, 846234000,
    846234900, 846235800, 846236700, 846237600, 846238500, 846239400,
    846240300, 846241200, 846242100, 846243000, 846243900, 846244800,
    846245700, 846246600, 846247500, 846248400, 846249300, 846250200,
    846251100, 846252000, 846252900, 846253800, 846254700, 846255600,
    846256500, 846257400, 846258300, 846259200, 846260100, 846261000,
    846261900, 846262800, 846263700, 846264600, 846265500, 846266400,
    846267300, 846268200, 846269100, 846270000, 846270900, 846271800,
    846272700, 846273600, 846274500, 846275400, 846276300, 846277200,
    846278100, 846279000, 846279900, 846280800, 846281700, 846282600,
    846283500, 846284400, 846285300, 846286200, 846287100, 846288000,
    846288900, 846289800, 846290700, 846291600, 846292500, 846293400,
    846294300, 846295200, 846296100, 846297000, 846297900, 846298800,
    846299700, 846300600, 846301500, 846302400, 846303300, 846304200,
    846305100, 846306000, 846306900, 846307800, 846308700, 846309600,
    846310500, 846311400, 846312300, 846313200, 846314100, 846315000,
    846315900, 846316800, 846317700, 846318600, 846319500, 846320400,
    846321300, 846322200, 846323100, 846324000, 846324900, 846325800,
    846326700, 846327600, 846328500, 846329400, 846330300, 846331200,
    846332100, 846333000, 846333900, 846334800, 846335700, 846336600,
    846337500, 846338400, 846339300, 846340200, 846341100, 846342000,
    846342900, 846343800, 846344700, 846345600, 846346500, 846347400,
    846348300, 846349200, 846350100, 846351000, 846351900, 846352800,
    846353700, 846354600, 846355500, 846356400, 846357300, 846358200,
    846359100, 846360000, 846360900, 846361800, 846362700, 846363600,
    846364500, 846365400, 846366300, 846367200, 846368100, 846369000,
    846369900, 846370800, 846371700, 846372600, 846373500, 846374400,
    846375300, 846376200, 846377100, 846378000, 846378900, 846379800,
    846380700, 846381600, 846382500, 846383400, 846384300, 846385200,
    846386100, 846387000, 846387900, 846388800, 846389700, 846390600,
    846391500, 846392400, 846393300, 846394200, 846395100, 846396000,
    846396900, 846397800, 846398700, 846399600, 846400500, 846401400,
    846402300, 846403200, 846404100, 846405000, 846405900, 846406800,
    846407700, 846408600, 846409500, 846410400, 846411300, 846412200,
    846413100, 846414000, 846414900, 846415800, 846416700, 846417600,
    846418500, 846419400, 846420300, 846421200, 846422100, 846423000,
    846423900, 846424800, 846425700, 846426600, 846427500, 846428400,
    846429300, 846430200, 846431100, 846432000, 846432900, 846433800,
    846434700, 846435600, 846436500, 846437400, 846438300, 846439200,
    846440100, 846441000, 846441900, 846442800, 846443700, 846444600,
    846445500, 846446400, 846447300, 846448200, 846449100, 846450000,
    846450900, 846451800, 846452700, 846453600, 846454500, 846455400,
    846456300, 846457200, 846458100, 846459000, 846459900, 846460800,
    846461700, 846462600, 846463500, 846464400, 846465300, 846466200,
    846467100, 846468000, 846468900, 846469800, 846470700, 846471600,
    846472500, 846473400, 846474300, 846475200, 846476100, 846477000,
    846477900, 846478800, 846479700, 846480600, 846481500, 846482400,
    846483300, 846484200, 846485100, 846486000, 846486900, 846487800,
    846488700, 846489600, 846490500, 846491400, 846492300, 846493200,
    846494100, 846495000, 846495900, 846496800, 846497700, 846498600,
    846499500, 846500400, 846501300, 846502200, 846503100, 846504000,
    846504900, 846505800, 846506700, 846507600, 846508500, 846509400,
    846510300, 846511200, 846512100, 846513000, 846513900, 846514800,
    846515700, 846516600, 846517500, 846518400, 846519300, 846520200,
    846521100, 846522000, 846522900, 846523800, 846524700, 846525600,
    846526500, 846527400, 846528300, 846529200, 846530100, 846531000,
    846531900, 846532800, 846533700, 846534600, 846535500, 846536400,
    846537300, 846538200, 846539100, 846540000, 846540900, 846541800,
    846542700, 846543600, 846544500, 846545400, 846546300, 846547200,
    846548100, 846549000, 846549900, 846550800, 846551700, 846552600,
    846553500, 846554400, 846555300, 846556200, 846557100, 846558000,
    846558900, 846559800, 846560700, 846561600, 846562500, 846563400,
    846564300, 846565200, 846566100, 846567000, 846567900, 846568800,
    846569700, 846570600, 846571500, 846572400, 846573300, 846574200,
    846575100, 846576000, 846576900, 846577800, 846578700, 846579600,
    846580500, 846581400, 846582300, 846583200, 846584100, 846585000,
    846585900, 846586800, 846587700, 846588600, 846589500, 846590400,
    846591300, 846592200, 846593100, 846594000, 846594900, 846595800,
    846596700, 846597600, 846598500, 846599400, 846600300, 846601200,
    846602100, 846603000, 846603900, 846604800, 846605700, 846606600,
    846607500, 846608400, 846609300, 846610200, 846611100, 846612000,
    846612900, 846613800, 846614700, 846615600, 846616500, 846617400,
    846618300, 846619200, 846620100, 846621000, 846621900, 846622800,
    846623700, 846624600, 846625500, 846626400, 846627300, 846628200,
    846629100, 846630000, 846630900, 846631800, 846632700, 846633600,
    846634500, 846635400, 846636300, 846637200, 846638100, 846639000,
    846639900, 846640800, 846641700, 846642600, 846643500, 846644400,
    846645300, 846646200, 846647100, 846648000, 846648900, 846649800,
    846650700, 846651600, 846652500, 846653400, 846654300, 846655200,
    846656100, 846657000, 846657900, 846658800, 846659700, 846660600,
    846661500, 846662400, 846663300, 846664200, 846665100, 846666000,
    846666900, 846667800, 846668700, 846669600, 846670500, 846671400,
    846672300, 846673200, 846674100, 846675000, 846675900, 846676800,
    846677700, 846678600, 846679500, 846680400, 846681300, 846682200,
    846683100, 846684000, 846684900, 846685800, 846686700, 846687600,
    846688500, 846689400, 846690300, 846691200, 846692100, 846693000,
    846693900, 846694800, 846695700, 846696600, 846697500, 846698400,
    846699300, 846700200, 846701100, 846702000, 846702900, 846703800,
    846704700, 846705600, 846706500, 846707400, 846708300, 846709200,
    846710100, 846711000, 846711900, 846712800, 846713700, 846714600,
    846715500, 846716400, 846717300, 846718200, 846719100, 846720000,
    846720900, 846721800, 846722700, 846723600, 846724500, 846725400,
    846726300, 846727200, 846728100, 846729000, 846729900, 846730800,
    846731700, 846732600, 846733500, 846734400, 846735300, 846736200,
    846737100, 846738000, 846738900, 846739800, 846740700, 846741600,
    846742500, 846743400, 846744300, 846745200, 846746100, 846747000,
    846747900, 846748800, 846749700, 846750600, 846751500, 846752400,
    846753300, 846754200, 846755100, 846756000, 846756900, 846757800,
    846758700, 846759600, 846760500, 846761400, 846762300, 846763200,
    846764100, 846765000, 846765900, 846766800, 846767700, 846768600,
    846769500, 846770400, 846771300, 846772200, 846773100, 846774000,
    846774900, 846775800, 846776700, 846777600, 846778500, 846779400,
    846780300, 846781200, 846782100, 846783000, 846783900, 846784800,
    846785700, 846786600, 846787500, 846788400, 846789300, 846790200,
    846791100, 846792000, 846792900, 846793800, 846794700, 846795600,
    846796500, 846797400, 846798300, 846799200, 846800100, 846801000,
    846801900, 846802800, 846803700, 846804600, 846805500, 846806400,
    846807300, 846808200, 846809100, 846810000, 846810900, 846811800,
    846812700, 846813600, 846814500, 846815400, 846816300, 846817200,
    846818100, 846819000, 846819900, 846820800, 846821700, 846822600,
    846823500, 846824400, 846825300, 846826200, 846827100, 846828000,
    846828900, 846829800, 846830700, 846831600, 846832500, 846833400,
    846834300, 846835200, 846836100, 846837000, 846837900, 846838800,
    846839700, 846840600, 846841500, 846842400, 846843300, 846844200,
    846845100, 846846000, 846846900, 846847800, 846848700, 846849600,
    846850500, 846851400, 846852300, 846853200, 846854100, 846855000,
    846855900, 846856800, 846857700, 846858600, 846859500, 846860400,
    846861300, 846862200, 846863100, 846864000, 846864900, 846865800,
    846866700, 846867600, 846868500, 846869400, 846870300, 846871200,
    846872100, 846873000, 846873900, 846874800, 846875700, 846876600,
    846877500, 846878400, 846879300, 846880200, 846881100, 846882000,
    846882900, 846883800, 846884700, 846885600, 846886500, 846887400,
    846888300, 846889200, 846890100, 846891000, 846891900, 846892800,
    846893700, 846894600, 846895500, 846896400, 846897300, 846898200,
    846899100, 846900000, 846900900, 846901800, 846902700, 846903600,
    846904500, 846905400, 846906300, 846907200, 846908100, 846909000,
    846909900, 846910800, 846911700, 846912600, 846913500, 846914400,
    846915300, 846916200, 846917100, 846918000, 846918900, 846919800,
    846920700, 846921600, 846922500, 846923400, 846924300, 846925200,
    846926100, 846927000, 846927900, 846928800, 846929700, 846930600,
    846931500, 846932400, 846933300, 846934200, 846935100, 846936000,
    846936900, 846937800, 846938700, 846939600, 846940500, 846941400,
    846942300, 846943200, 846944100, 846945000, 846945900, 846946800,
    846947700, 846948600, 846949500, 846950400, 846951300, 846952200,
    846953100, 846954000, 846954900, 846955800, 846956700, 846957600,
    846958500, 846959400, 846960300, 846961200, 846962100, 846963000,
    846963900, 846964800, 846965700, 846966600, 846967500, 846968400,
    846969300, 846970200, 846971100, 846972000, 846972900, 846973800,
    846974700, 846975600, 846976500, 846977400, 846978300, 846979200,
    846980100, 846981000, 846981900, 846982800, 846983700, 846984600,
    846985500, 846986400, 846987300, 846988200, 846989100, 846990000,
    846990900, 846991800, 846992700, 846993600, 846994500, 846995400,
    846996300, 846997200, 846998100, 846999000, 846999900, 847000800,
    847001700, 847002600, 847003500, 847004400, 847005300, 847006200,
    847007100, 847008000, 847008900, 847009800, 847010700, 847011600,
    847012500, 847013400, 847014300, 847015200, 847016100, 847017000,
    847017900, 847018800, 847019700, 847020600, 847021500, 847022400,
    847023300, 847024200, 847025100, 847026000, 847026900, 847027800,
    847028700, 847029600, 847030500, 847031400, 847032300, 847033200,
    847034100, 847035000, 847035900, 847036800, 847037700, 847038600,
    847039500, 847040400, 847041300, 847042200, 847043100, 847044000,
    847044900, 847045800, 847046700, 847047600, 847048500, 847049400,
    847050300, 847051200, 847052100, 847053000, 847053900, 847054800,
    847055700, 847056600, 847057500, 847058400, 847059300, 847060200,
    847061100, 847062000, 847062900, 847063800, 847064700, 847065600,
    847066500, 847067400, 847068300, 847069200, 847070100, 847071000,
    847071900, 847072800, 847073700, 847074600, 847075500, 847076400,
    847077300, 847078200, 847079100, 847080000, 847080900, 847081800,
    847082700, 847083600, 847084500, 847085400, 847086300, 847087200,
    847088100, 847089000, 847089900, 847090800, 847091700, 847092600,
    847093500, 847094400, 847095300, 847096200, 847097100, 847098000,
    847098900, 847099800, 847100700, 847101600, 847102500, 847103400,
    847104300, 847105200, 847106100, 847107000, 847107900, 847108800,
    847109700, 847110600, 847111500, 847112400, 847113300, 847114200,
    847115100, 847116000, 847116900, 847117800, 847118700, 847119600,
    847120500, 847121400, 847122300, 847123200, 847124100, 847125000,
    847125900, 847126800, 847127700, 847128600, 847129500, 847130400,
    847131300, 847132200, 847133100, 847134000, 847134900, 847135800,
    847136700, 847137600, 847138500, 847139400, 847140300, 847141200,
    847142100, 847143000, 847143900, 847144800, 847145700, 847146600,
    847147500, 847148400, 847149300, 847150200, 847151100, 847152000,
    847152900, 847153800, 847154700, 847155600, 847156500, 847157400,
    847158300, 847159200, 847160100, 847161000, 847161900, 847162800,
    847163700, 847164600, 847165500, 847166400, 847167300, 847168200,
    847169100, 847170000, 847170900, 847171800, 847172700, 847173600,
    847174500, 847175400, 847176300, 847177200, 847178100, 847179000,
    847179900, 847180800, 847181700, 847182600, 847183500, 847184400,
    847185300, 847186200, 847187100, 847188000, 847188900, 847189800,
    847190700, 847191600, 847192500, 847193400, 847194300, 847195200,
    847196100, 847197000, 847197900, 847198800, 847199700, 847200600,
    847201500, 847202400, 847203300, 847204200, 847205100, 847206000,
    847206900, 847207800, 847208700, 847209600, 847210500, 847211400,
    847212300, 847213200, 847214100, 847215000, 847215900, 847216800,
    847217700, 847218600, 847219500, 847220400, 847221300, 847222200,
    847223100, 847224000, 847224900, 847225800, 847226700, 847227600,
    847228500, 847229400, 847230300, 847231200, 847232100, 847233000,
    847233900, 847234800, 847235700, 847236600, 847237500, 847238400,
    847239300, 847240200, 847241100, 847242000, 847242900, 847243800,
    847244700, 847245600, 847246500, 847247400, 847248300, 847249200,
    847250100, 847251000, 847251900, 847252800, 847253700, 847254600,
    847255500, 847256400, 847257300, 847258200, 847259100, 847260000,
    847260900, 847261800, 847262700, 847263600, 847264500, 847265400,
    847266300, 847267200, 847268100, 847269000, 847269900, 847270800,
    847271700, 847272600, 847273500, 847274400, 847275300, 847276200,
    847277100, 847278000, 847278900, 847279800, 847280700, 847281600,
    847282500, 847283400, 847284300, 847285200, 847286100, 847287000,
    847287900, 847288800, 847289700, 847290600, 847291500, 847292400,
    847293300, 847294200, 847295100, 847296000, 847296900, 847297800,
    847298700, 847299600, 847300500, 847301400, 847302300, 847303200,
    847304100, 847305000, 847305900, 847306800, 847307700, 847308600,
    847309500, 847310400, 847311300, 847312200, 847313100, 847314000,
    847314900, 847315800, 847316700, 847317600, 847318500, 847319400,
    847320300, 847321200, 847322100, 847323000, 847323900, 847324800,
    847325700, 847326600, 847327500, 847328400, 847329300, 847330200,
    847331100, 847332000, 847332900, 847333800, 847334700, 847335600,
    847336500, 847337400, 847338300, 847339200, 847340100, 847341000,
    847341900, 847342800, 847343700, 847344600, 847345500, 847346400,
    847347300, 847348200, 847349100, 847350000, 847350900, 847351800,
    847352700, 847353600, 847354500, 847355400, 847356300, 847357200,
    847358100, 847359000, 847359900, 847360800, 847361700, 847362600,
    847363500, 847364400, 847365300, 847366200, 847367100, 847368000,
    847368900, 847369800, 847370700, 847371600, 847372500, 847373400,
    847374300, 847375200, 847376100, 847377000, 847377900, 847378800,
    847379700, 847380600, 847381500, 847382400, 847383300, 847384200,
    847385100, 847386000, 847386900, 847387800, 847388700, 847389600,
    847390500, 847391400, 847392300, 847393200, 847394100, 847395000,
    847395900, 847396800, 847397700, 847398600, 847399500, 847400400,
    847401300, 847402200, 847403100, 847404000, 847404900, 847405800,
    847406700, 847407600, 847408500, 847409400, 847410300, 847411200,
    847412100, 847414800, 847415700, 847416600, 847417500, 847418400,
    847419300, 847420200, 847421100, 847422000, 847422900, 847423800,
    847424700, 847425600, 847426500, 847427400, 847428300, 847429200,
    847430100, 847431000, 847431900, 847432800, 847433700, 847434600,
    847435500, 847436400, 847437300, 847438200, 847439100, 847440000,
    847440900, 847441800, 847442700, 847443600, 847444500, 847445400,
    847446300, 847447200, 847448100, 847449000, 847449900, 847450800,
    847451700, 847452600, 847453500, 847454400, 847455300, 847456200,
    847457100, 847458000, 847458900, 847459800, 847460700, 847461600,
    847462500, 847463400, 847464300, 847465200, 847466100, 847467000,
    847467900, 847468800, 847469700, 847470600, 847471500, 847472400,
    847473300, 847474200, 847475100, 847476000, 847476900, 847477800,
    847478700, 847479600, 847480500, 847481400, 847482300, 847483200,
    847484100, 847485000, 847485900, 847486800, 847487700, 847488600,
    847489500, 847490400, 847491300, 847492200, 847493100, 847494000,
    847494900, 847495800, 847496700, 847497600, 847498500, 847499400,
    847500300, 847501200, 847502100, 847503000, 847503900, 847504800,
    847505700, 847506600, 847507500, 847508400, 847509300, 847510200,
    847511100, 847512000, 847512900, 847513800, 847514700, 847515600,
    847516500, 847517400, 847518300, 847519200, 847520100, 847521000,
    847521900, 847522800, 847523700, 847524600, 847525500, 847526400,
    847527300, 847528200, 847529100, 847530000, 847530900, 847531800,
    847532700, 847533600, 847534500, 847535400, 847536300, 847537200,
    847538100, 847539000, 847539900, 847540800, 847541700, 847542600,
    847543500, 847544400, 847545300, 847546200, 847547100, 847548000,
    847548900, 847549800, 847550700, 847551600, 847552500, 847553400,
    847554300, 847555200, 847556100, 847557000, 847557900, 847558800,
    847559700, 847560600, 847561500, 847562400, 847563300, 847564200,
    847565100, 847566000, 847566900, 847567800, 847568700, 847569600,
    847570500, 847571400, 847572300, 847573200, 847574100, 847575000,
    847575900, 847576800, 847577700, 847578600, 847579500, 847580400,
    847581300, 847582200, 847583100, 847584000, 847584900, 847585800,
    847586700, 847587600, 847588500, 847589400, 847590300, 847591200,
    847592100, 847593000, 847593900, 847594800, 847595700, 847596600,
    847597500, 847598400, 847599300, 847600200, 847601100, 847602000,
    847602900, 847603800, 847604700, 847605600, 847606500, 847607400,
    847608300, 847609200, 847610100, 847611000, 847611900, 847612800,
    847613700, 847614600, 847615500, 847616400, 847617300, 847618200,
    847619100, 847620000, 847620900, 847621800, 847622700, 847623600,
    847624500, 847625400, 847626300, 847627200, 847628100, 847629000,
    847629900, 847630800, 847631700, 847632600, 847633500, 847634400,
    847635300, 847636200, 847637100, 847638000, 847638900, 847639800,
    847640700, 847641600, 847642500, 847643400, 847644300, 847645200,
    847646100, 847647000, 847647900, 847648800, 847649700, 847650600,
    847651500, 847652400, 847653300, 847654200, 847655100, 847656000,
    847656900, 847657800, 847658700, 847659600, 847660500, 847661400,
    847662300, 847663200, 847664100, 847665000, 847665900, 847666800,
    847667700, 847668600, 847669500, 847670400, 847671300, 847672200,
    847673100, 847674000, 847674900, 847675800, 847676700, 847677600,
    847678500, 847679400, 847680300, 847681200, 847682100, 847683000,
    847683900, 847684800, 847685700, 847686600, 847687500, 847688400,
    847689300, 847690200, 847691100, 847692000, 847692900, 847693800,
    847694700, 847695600, 847696500, 847697400, 847698300, 847699200,
    847700100, 847701000, 847701900, 847702800, 847703700, 847704600,
    847705500, 847706400, 847707300, 847708200, 847709100, 847710000,
    847710900, 847711800, 847712700, 847713600, 847714500, 847715400,
    847716300, 847717200, 847718100, 847719000, 847719900, 847720800,
    847721700, 847722600, 847723500, 847724400, 847725300, 847726200,
    847727100, 847728000, 847728900, 847729800, 847730700, 847731600,
    847732500, 847733400, 847734300, 847735200, 847736100, 847737000,
    847737900, 847738800, 847739700, 847740600, 847741500, 847742400,
    847743300, 847744200, 847745100, 847746000, 847746900, 847747800,
    847748700, 847749600, 847750500, 847751400, 847752300, 847753200,
    847754100, 847755000, 847755900, 847756800, 847757700, 847758600,
    847759500, 847760400, 847761300, 847762200, 847763100, 847764000,
    847764900, 847765800, 847766700, 847767600, 847768500, 847769400,
    847770300, 847771200, 847772100, 847773000, 847773900, 847774800,
    847775700, 847776600, 847777500, 847778400, 847779300, 847780200,
    847781100, 847782000, 847782900, 847783800, 847784700, 847785600,
    847786500, 847787400, 847788300, 847789200, 847790100, 847791000,
    847791900, 847792800, 847793700, 847794600, 847795500, 847796400,
    847797300, 847798200, 847799100, 847800000, 847800900, 847801800,
    847802700, 847803600, 847804500, 847805400, 847806300, 847807200,
    847808100, 847809000, 847809900, 847810800, 847811700, 847812600,
    847813500, 847814400, 847815300, 847816200, 847817100, 847818000,
    847818900, 847819800, 847820700, 847821600, 847822500, 847823400,
    847824300, 847825200, 847826100, 847827000, 847827900, 847828800,
    847829700, 847830600, 847831500, 847832400, 847833300, 847834200,
    847835100, 847836000, 847836900, 847837800, 847838700, 847839600,
    847840500, 847841400, 847842300, 847843200, 847844100, 847845000,
    847845900, 847846800, 847847700, 847848600, 847849500, 847850400,
    847851300, 847852200, 847853100, 847854000, 847854900, 847855800,
    847856700, 847857600, 847858500, 847859400, 847860300, 847861200,
    847862100, 847863000, 847863900, 847864800, 847865700, 847866600,
    847867500, 847868400, 847869300, 847870200, 847871100, 847872000,
    847872900, 847873800, 847874700, 847875600, 847876500, 847877400,
    847878300, 847879200, 847880100, 847881000, 847881900, 847882800,
    847883700, 847884600, 847885500, 847886400, 847887300, 847888200,
    847889100, 847890000, 847890900, 847891800, 847892700, 847893600,
    847894500, 847895400, 847896300, 847897200, 847898100, 847899000,
    847899900, 847900800, 847901700, 847902600, 847903500, 847904400,
    847905300, 847906200, 847907100, 847908000, 847908900, 847909800,
    847910700, 847911600, 847912500, 847913400, 847914300, 847915200,
    847916100, 847917000, 847917900, 847918800, 847919700, 847920600,
    847921500, 847922400, 847923300, 847924200, 847925100, 847926000,
    847926900, 847927800, 847928700, 847929600, 847930500, 847931400,
    847932300, 847933200, 847934100, 847935000, 847935900, 847936800,
    847937700, 847938600, 847939500, 847940400, 847941300, 847942200,
    847943100, 847944000, 847944900, 847945800, 847946700, 847947600,
    847948500, 847949400, 847950300, 847951200, 847952100, 847953000,
    847953900, 847954800, 847955700, 847956600, 847957500, 847958400,
    847959300, 847960200, 847961100, 847962000, 847962900, 847963800,
    847964700, 847965600, 847966500, 847967400, 847968300, 847969200,
    847970100, 847971000, 847971900, 847972800, 847973700, 847974600,
    847975500, 847976400, 847977300, 847978200, 847979100, 847980000,
    847980900, 847981800, 847982700, 847983600, 847984500, 847985400,
    847986300, 847987200, 847988100, 847989000, 847989900, 847990800,
    847991700, 847992600, 847993500, 847994400, 847995300, 847996200,
    847997100, 847998000, 847998900, 847999800, 848000700, 848001600,
    848002500, 848003400, 848004300, 848005200, 848006100, 848007000,
    848007900, 848008800, 848009700, 848010600, 848011500, 848012400,
    848013300, 848014200, 848015100, 848016000, 848016900, 848017800,
    848018700, 848019600, 848020500, 848021400, 848022300, 848023200,
    848024100, 848025000, 848025900, 848026800, 848027700, 848028600,
    848029500, 848030400, 848031300, 848032200, 848033100, 848034000,
    848034900, 848035800, 848036700, 848037600, 848038500, 848039400,
    848040300, 848041200, 848042100, 848043000, 848043900, 848044800,
    848045700, 848046600, 848047500, 848048400, 848049300, 848050200,
    848051100, 848052000, 848052900, 848053800, 848054700, 848055600,
    848056500, 848057400, 848058300, 848059200, 848060100, 848061000,
    848061900, 848062800, 848063700, 848064600, 848065500, 848066400,
    848067300, 848068200, 848069100, 848070000, 848070900, 848071800,
    848072700, 848073600, 848074500, 848075400, 848076300, 848077200,
    848078100, 848079000, 848079900, 848080800, 848081700, 848082600,
    848083500, 848084400, 848085300, 848086200, 848087100, 848088000,
    848088900, 848089800, 848090700, 848091600, 848092500, 848093400,
    848094300, 848095200, 848096100, 848097000, 848097900, 848098800,
    848099700, 848100600, 848101500, 848102400, 848103300, 848104200,
    848105100, 848106000, 848106900, 848107800, 848108700, 848109600,
    848110500, 848111400, 848112300, 848113200, 848114100, 848115000,
    848115900, 848116800, 848117700, 848118600, 848119500, 848120400,
    848121300, 848122200, 848123100, 848124000, 848124900, 848125800,
    848126700, 848127600, 848128500, 848129400, 848130300, 848131200,
    848132100, 848133000, 848133900, 848134800, 848135700, 848136600,
    848137500, 848138400, 848139300, 848140200, 848141100, 848142000,
    848142900, 848143800, 848144700, 848145600, 848146500, 848147400,
    848148300, 848149200, 848150100, 848151000, 848151900, 848152800,
    848153700, 848154600, 848155500, 848156400, 848157300, 848158200,
    848159100, 848160000, 848160900, 848161800, 848162700, 848163600,
    848164500, 848165400, 848166300, 848167200, 848168100, 848169000,
    848169900, 848170800, 848171700, 848172600, 848173500, 848174400,
    848175300, 848176200, 848177100, 848178000, 848178900, 848179800,
    848180700, 848181600, 848182500, 848183400, 848184300, 848185200,
    848186100, 848187000, 848187900, 848188800, 848189700, 848190600,
    848191500, 848192400, 848193300, 848194200, 848195100, 848196000,
    848196900, 848197800, 848198700, 848199600, 848200500, 848201400,
    848202300, 848203200, 848204100, 848205000, 848205900, 848206800,
    848207700, 848208600, 848209500, 848210400, 848211300, 848212200,
    848213100, 848214000, 848214900, 848215800, 848216700, 848217600,
    848218500, 848219400, 848220300, 848221200, 848222100, 848223000,
    848223900, 848224800, 848225700, 848226600, 848227500, 848228400,
    848229300, 848230200, 848231100, 848232000, 848232900, 848233800,
    848234700, 848235600, 848236500, 848237400, 848238300, 848239200,
    848240100, 848241000, 848241900, 848242800, 848243700, 848244600,
    848245500, 848246400, 848247300, 848248200, 848249100, 848250000,
    848250900, 848251800, 848252700, 848253600, 848254500, 848255400,
    848256300, 848257200, 848258100, 848259000, 848259900, 848260800,
    848261700, 848262600, 848263500, 848264400, 848265300, 848266200,
    848267100, 848268000, 848268900, 848269800, 848270700, 848271600,
    848272500, 848273400, 848274300, 848275200, 848276100, 848277000,
    848277900, 848278800, 848279700, 848280600, 848281500, 848282400,
    848283300, 848284200, 848285100, 848286000, 848286900, 848287800,
    848288700, 848289600, 848290500, 848291400, 848292300, 848293200,
    848294100, 848295000, 848295900, 848296800, 848297700, 848298600,
    848299500, 848300400, 848301300, 848302200, 848303100, 848304000,
    848304900, 848305800, 848306700, 848307600, 848308500, 848309400,
    848310300, 848311200, 848312100, 848313000, 848313900, 848314800,
    848315700, 848316600, 848317500, 848318400, 848319300, 848320200,
    848321100, 848322000, 848322900, 848323800, 848324700, 848325600,
    848326500, 848327400, 848328300, 848329200, 848330100, 848331000,
    848331900, 848332800, 848333700, 848334600, 848335500, 848336400,
    848337300, 848338200, 848339100, 848340000, 848340900, 848341800,
    848342700, 848343600, 848344500, 848345400, 848346300, 848347200,
    848348100, 848349000, 848349900, 848350800, 848351700, 848352600,
    848353500, 848354400, 848355300, 848356200, 848357100, 848358000,
    848358900, 848359800, 848360700, 848361600, 848362500, 848363400,
    848364300, 848365200, 848366100, 848367000, 848367900, 848368800,
    848369700, 848370600, 848371500, 848372400, 848373300, 848374200,
    848375100, 848376000, 848376900, 848377800, 848378700, 848379600,
    848380500, 848381400, 848382300, 848383200, 848384100, 848385000,
    848385900, 848386800, 848387700, 848388600, 848389500, 848390400,
    848391300, 848392200, 848393100, 848394000, 848394900, 848395800,
    848396700, 848397600, 848398500, 848399400, 848400300, 848401200,
    848402100, 848403000, 848403900, 848404800, 848405700, 848406600,
    848407500, 848408400, 848409300, 848410200, 848411100, 848412000,
    848412900, 848413800, 848414700, 848415600, 848416500, 848417400,
    848418300, 848419200, 848420100, 848421000, 848421900, 848422800,
    848423700, 848424600, 848425500, 848426400, 848427300, 848428200,
    848429100, 848430000, 848430900, 848431800, 848432700, 848433600,
    848434500, 848435400, 848436300, 848437200, 848438100, 848439000,
    848439900, 848440800, 848441700, 848442600, 848443500, 848444400,
    848445300, 848446200, 848447100, 848448000, 848448900, 848449800,
    848450700, 848451600, 848452500, 848453400, 848454300, 848455200,
    848456100, 848457000, 848457900, 848458800, 848459700, 848460600,
    848461500, 848462400, 848463300, 848464200, 848465100, 848466000,
    848466900, 848467800, 848468700, 848469600, 848470500, 848471400,
    848472300, 848473200, 848474100, 848475000, 848475900, 848476800,
    848477700, 848478600, 848479500, 848480400, 848481300, 848482200,
    848483100, 848484000, 848484900, 848485800, 848486700, 848487600,
    848488500, 848489400, 848490300, 848491200, 848492100, 848493000,
    848493900, 848494800, 848495700, 848496600, 848497500, 848498400,
    848499300, 848500200, 848501100, 848502000, 848502900, 848503800,
    848504700, 848505600, 848506500, 848507400, 848508300, 848509200,
    848510100, 848511000, 848511900, 848512800, 848513700, 848514600,
    848515500, 848516400, 848517300, 848518200, 848519100, 848520000,
    848520900, 848521800, 848522700, 848523600, 848524500, 848525400,
    848526300, 848527200, 848528100, 848529000, 848529900, 848530800,
    848531700, 848532600, 848533500, 848534400, 848535300, 848536200,
    848537100, 848538000, 848538900, 848539800, 848540700, 848541600,
    848542500, 848543400, 848544300, 848545200, 848546100, 848547000,
    848547900, 848548800, 848549700, 848550600, 848551500, 848552400,
    848553300, 848554200, 848555100, 848556000, 848556900, 848557800,
    848558700, 848559600, 848560500, 848561400, 848562300, 848563200,
    848564100, 848565000, 848565900, 848566800, 848567700, 848568600,
    848569500, 848570400, 848571300, 848572200, 848573100, 848574000,
    848574900, 848575800, 848576700, 848577600, 848578500, 848579400,
    848580300, 848581200, 848582100, 848583000, 848583900, 848584800,
    848585700, 848586600, 848587500, 848588400, 848589300, 848590200,
    848591100, 848592000, 848592900, 848593800, 848594700, 848595600,
    848596500, 848597400, 848598300, 848599200, 848600100, 848601000,
    848601900, 848602800, 848603700, 848604600, 848605500, 848606400,
    848607300, 848608200, 848609100, 848610000, 848610900, 848611800,
    848612700, 848613600, 848614500, 848615400, 848616300, 848617200,
    848618100, 848619000, 848619900, 848620800, 848621700, 848622600,
    848623500, 848624400, 848625300, 848626200, 848627100, 848628000,
    848628900, 848629800, 848630700, 848631600, 848632500, 848633400,
    848634300, 848635200, 848636100, 848637000, 848637900, 848638800,
    848639700, 848640600, 848641500, 848642400, 848643300, 848644200,
    848645100, 848646000, 848646900, 848647800, 848648700, 848649600,
    848650500, 848651400, 848652300, 848653200, 848654100, 848655000,
    848655900, 848656800, 848657700, 848658600, 848659500, 848660400,
    848661300, 848662200, 848663100, 848664000, 848664900, 848665800,
    848666700, 848667600, 848668500, 848669400, 848670300, 848671200,
    848672100, 848673000, 848673900, 848674800, 848675700, 848676600,
    848677500, 848678400, 848679300, 848680200, 848681100, 848682000,
    848682900, 848683800, 848684700, 848685600, 848686500, 848687400,
    848688300, 848689200, 848690100, 848691000, 848691900, 848692800,
    848693700, 848694600, 848695500, 848696400, 848697300, 848698200,
    848699100, 848700000, 848700900, 848701800, 848702700, 848703600,
    848704500, 848705400, 848706300, 848707200, 848708100, 848709000,
    848709900, 848710800, 848711700, 848712600, 848713500, 848714400,
    848715300, 848716200, 848717100, 848718000, 848718900, 848719800,
    848720700, 848721600, 848722500, 848723400, 848724300, 848725200,
    848726100, 848727000, 848727900, 848728800, 848729700, 848730600,
    848731500, 848732400, 848733300, 848734200, 848735100, 848736000,
    848736900, 848737800, 848738700, 848739600, 848740500, 848741400,
    848742300, 848743200, 848744100, 848745000, 848745900, 848746800,
    848747700, 848748600, 848749500, 848750400, 848751300, 848752200,
    848753100, 848754000, 848754900, 848755800, 848756700, 848757600,
    848758500, 848759400, 848760300, 848761200, 848762100, 848763000,
    848763900, 848764800, 848765700, 848766600, 848767500, 848768400,
    848769300, 848770200, 848771100, 848772000, 848772900, 848773800,
    848774700, 848775600, 848776500, 848777400, 848778300, 848779200,
    848780100, 848781000, 848781900, 848782800, 848783700, 848784600,
    848785500, 848786400, 848787300, 848788200, 848789100, 848790000,
    848790900, 848791800, 848792700, 848793600, 848794500, 848795400,
    848796300, 848797200, 848798100, 848799000, 848799900, 848800800,
    848801700, 848802600, 848803500, 848804400, 848805300, 848806200,
    848807100, 848808000, 848808900, 848809800, 848810700, 848811600,
    848812500, 848813400, 848814300, 848815200, 848816100, 848817000,
    848817900, 848818800, 848819700, 848820600, 848821500, 848822400,
    848823300, 848824200, 848825100, 848826000, 848826900, 848827800,
    848828700, 848829600, 848830500, 848831400, 848832300, 848833200,
    848834100, 848835000, 848835900, 848836800, 848837700, 848838600,
    848839500, 848840400, 848841300, 848842200, 848843100, 848844000,
    848844900, 848845800, 848846700, 848847600, 848848500, 848849400,
    848850300, 848851200, 848852100, 848853000, 848853900, 848854800,
    848855700, 848856600, 848857500, 848858400, 848859300, 848860200,
    848861100, 848862000, 848862900, 848863800, 848864700, 848865600,
    848866500, 848867400, 848868300, 848869200, 848870100, 848871000,
    848871900, 848872800, 848873700, 848874600, 848875500, 848876400,
    848877300, 848878200, 848879100, 848880000, 848880900, 848881800,
    848882700, 848883600, 848884500, 848885400, 848886300, 848887200,
    848888100, 848889000, 848889900, 848890800, 848891700, 848892600,
    848893500, 848894400, 848895300, 848896200, 848897100, 848898000,
    848898900, 848899800, 848900700, 848901600, 848902500, 848903400,
    848904300, 848905200, 848906100, 848907000, 848907900, 848908800,
    848909700, 848910600, 848911500, 848912400, 848913300, 848914200,
    848915100, 848916000, 848916900, 848917800, 848918700, 848919600,
    848920500, 848921400, 848922300, 848923200, 848924100, 848925000,
    848925900, 848926800, 848927700, 848928600, 848929500, 848930400,
    848931300, 848932200, 848933100, 848934000, 848934900, 848935800,
    848936700, 848937600, 848938500, 848939400, 848940300, 848941200,
    848942100, 848943000, 848943900, 848944800, 848945700, 848946600,
    848947500, 848948400, 848949300, 848950200, 848951100, 848952000,
    848952900, 848953800, 848954700, 848955600, 848956500, 848957400,
    848958300, 848959200, 848960100, 848961000, 848961900, 848962800,
    848963700, 848964600, 848965500, 848966400, 848967300, 848968200,
    848969100, 848970000, 848970900, 848971800, 848972700, 848973600,
    848974500, 848975400, 848976300, 848977200, 848978100, 848979000,
    848979900, 848980800, 848981700, 848982600, 848983500, 848984400,
    848985300, 848986200, 848987100, 848988000, 848988900, 848989800,
    848990700, 848991600, 848992500, 848993400, 848994300, 848995200,
    848996100, 848997000, 848997900, 848998800, 848999700, 849000600,
    849001500, 849002400, 849003300, 849004200, 849005100, 849006000,
    849006900, 849007800, 849008700, 849009600, 849010500, 849011400,
    849012300, 849013200, 849014100, 849015000, 849015900, 849016800,
    849017700, 849018600, 849019500, 849020400, 849021300, 849022200,
    849023100, 849024000, 849024900, 849025800, 849026700, 849027600,
    849028500, 849029400, 849030300, 849031200, 849032100, 849033000,
    849033900, 849034800, 849035700, 849036600, 849037500, 849038400,
    849039300, 849040200, 849041100, 849042000, 849042900, 849043800,
    849044700, 849045600, 849046500, 849047400, 849048300, 849049200,
    849050100, 849051000, 849051900, 849052800, 849053700, 849054600,
    849055500, 849056400, 849057300, 849058200, 849059100, 849060000,
    849060900, 849061800, 849062700, 849063600, 849064500, 849065400,
    849066300, 849067200, 849068100, 849069000, 849069900, 849070800,
    849071700, 849072600, 849073500, 849074400, 849075300, 849076200,
    849077100, 849078000, 849078900, 849079800, 849080700, 849081600,
    849082500, 849083400, 849084300, 849085200, 849086100, 849087000,
    849087900, 849088800, 849089700, 849090600, 849091500, 849092400,
    849093300, 849094200, 849095100, 849096000, 849096900, 849097800,
    849098700, 849099600, 849100500, 849101400, 849102300, 849103200,
    849104100, 849105000, 849105900, 849106800, 849107700, 849108600,
    849109500, 849110400, 849111300, 849112200, 849113100, 849114000,
    849114900, 849115800, 849116700, 849117600, 849118500, 849119400,
    849120300, 849121200, 849122100, 849123000, 849123900, 849124800,
    849125700, 849126600, 849127500, 849128400, 849129300, 849130200,
    849131100, 849132000, 849132900, 849133800, 849134700, 849135600,
    849136500, 849137400, 849138300, 849139200, 849140100, 849141000,
    849141900, 849142800, 849143700, 849144600, 849145500, 849146400,
    849147300, 849148200, 849149100, 849150000, 849150900, 849151800,
    849152700, 849153600, 849154500, 849155400, 849156300, 849157200,
    849158100, 849159000, 849159900, 849160800, 849161700, 849162600,
    849163500, 849164400, 849165300, 849166200, 849167100, 849168000,
    849168900, 849169800, 849170700, 849171600, 849172500, 849173400,
    849174300, 849175200, 849176100, 849177000, 849177900, 849178800,
    849179700, 849180600, 849181500, 849182400, 849183300, 849184200,
    849185100, 849186000, 849186900, 849187800, 849188700, 849189600,
    849190500, 849191400, 849192300, 849193200, 849194100, 849195000,
    849195900, 849196800, 849197700, 849198600, 849199500, 849200400,
    849201300, 849202200, 849203100, 849204000, 849204900, 849205800,
    849206700, 849207600, 849208500, 849209400, 849210300, 849211200,
    849212100, 849213000, 849213900, 849214800, 849215700, 849216600,
    849217500, 849218400, 849219300, 849220200, 849221100, 849222000,
    849222900, 849223800, 849224700, 849225600, 849226500, 849227400,
    849228300, 849229200, 849230100, 849231000, 849231900, 849232800,
    849233700, 849234600, 849235500, 849236400, 849237300, 849238200,
    849239100, 849240000, 849240900, 849241800, 849242700, 849243600,
    849244500, 849245400, 849246300, 849247200, 849248100, 849249000,
    849249900, 849250800, 849251700, 849252600, 849253500, 849254400,
    849255300, 849256200, 849257100, 849258000, 849258900, 849259800,
    849260700, 849261600, 849262500, 849263400, 849264300, 849265200,
    849266100, 849267000, 849267900, 849268800, 849269700, 849270600,
    849271500, 849272400, 849273300, 849274200, 849275100, 849276000,
    849276900, 849277800, 849278700, 849279600, 849280500, 849281400,
    849282300, 849283200, 849284100, 849285000, 849285900, 849286800,
    849287700, 849288600, 849289500, 849290400, 849291300, 849292200,
    849293100, 849294000, 849294900, 849295800, 849296700, 849297600,
    849298500, 849299400, 849300300, 849301200, 849302100, 849303000,
    849303900, 849304800, 849305700, 849306600, 849307500, 849308400,
    849309300, 849310200, 849311100, 849312000, 849312900, 849313800,
    849314700, 849315600, 849316500, 849317400, 849318300, 849319200,
    849320100, 849321000, 849321900, 849322800, 849323700, 849324600,
    849325500, 849326400, 849327300, 849328200, 849329100, 849330000,
    849330900, 849331800, 849332700, 849333600, 849334500, 849335400,
    849336300, 849337200, 849338100, 849339000, 849339900, 849340800,
    849341700, 849342600, 849343500, 849344400, 849345300, 849346200,
    849347100, 849348000, 849348900, 849349800, 849350700, 849351600,
    849352500, 849353400, 849354300, 849355200, 849356100, 849357000,
    849357900, 849358800, 849359700, 849360600, 849361500, 849362400,
    849363300, 849364200, 849365100, 849366000, 849366900, 849367800,
    849368700, 849369600, 849370500, 849371400, 849372300, 849373200,
    849374100, 849375000, 849375900, 849376800, 849377700, 849378600,
    849379500, 849380400, 849381300, 849382200, 849383100, 849384000,
    849384900, 849385800, 849386700, 849387600, 849388500, 849389400,
    849390300, 849391200, 849392100, 849393000, 849393900, 849394800,
    849395700, 849396600, 849397500, 849398400, 849399300, 849400200,
    849401100, 849402000, 849402900, 849403800, 849404700, 849405600,
    849406500, 849407400, 849408300, 849409200, 849410100, 849411000,
    849411900, 849412800, 849413700, 849414600, 849415500, 849416400,
    849417300, 849418200, 849419100, 849420000, 849420900, 849421800,
    849422700, 849423600, 849424500, 849425400, 849426300, 849427200,
    849428100, 849429000, 849429900, 849430800, 849431700, 849432600,
    849433500, 849434400, 849435300, 849436200, 849437100, 849438000,
    849438900, 849439800, 849440700, 849441600, 849442500, 849443400,
    849444300, 849445200, 849446100, 849447000, 849447900, 849448800,
    849449700, 849450600, 849451500, 849452400, 849453300, 849454200,
    849455100, 849456000, 849456900, 849457800, 849458700, 849459600,
    849460500, 849461400, 849462300, 849463200, 849464100, 849465000,
    849465900, 849466800, 849467700, 849468600, 849469500, 849470400,
    849471300, 849472200, 849473100, 849474000, 849474900, 849475800,
    849476700, 849477600, 849478500, 849479400, 849480300, 849481200,
    849482100, 849483000, 849483900, 849484800, 849485700, 849486600,
    849487500, 849488400, 849489300, 849490200, 849491100, 849492000,
    849492900, 849493800, 849494700, 849495600, 849496500, 849497400,
    849498300, 849499200, 849500100, 849501000, 849501900, 849502800,
    849503700, 849504600, 849505500, 849506400, 849507300, 849508200,
    849509100, 849510000, 849510900, 849511800, 849512700, 849513600,
    849514500, 849515400, 849516300, 849517200, 849518100, 849519000,
    849519900, 849520800, 849521700, 849522600, 849523500, 849524400,
    849525300, 849526200, 849527100, 849528000, 849528900, 849529800,
    849530700, 849531600, 849532500, 849533400, 849534300, 849535200,
    849536100, 849537000, 849537900, 849538800, 849539700, 849540600,
    849541500, 849542400, 849543300, 849544200, 849545100, 849546000,
    849546900, 849547800, 849548700, 849549600, 849550500, 849551400,
    849552300, 849553200, 849554100, 849555000, 849555900, 849556800,
    849557700, 849558600, 849559500, 849560400, 849561300, 849562200,
    849563100, 849564000, 849564900, 849565800, 849566700, 849567600,
    849568500, 849569400, 849570300, 849571200, 849572100, 849573000,
    849573900, 849574800, 849575700, 849576600, 849577500, 849578400,
    849579300, 849580200, 849581100, 849582000, 849582900, 849583800,
    849584700, 849585600, 849586500, 849587400, 849588300, 849589200,
    849590100, 849591000, 849591900, 849592800, 849593700, 849594600,
    849595500, 849596400, 849597300, 849598200, 849599100, 849600000,
    849600900, 849601800, 849602700, 849603600, 849604500, 849605400,
    849606300, 849607200, 849608100, 849609000, 849609900, 849610800,
    849611700, 849612600, 849613500, 849614400, 849615300, 849616200,
    849617100, 849618000, 849618900, 849619800, 849620700, 849621600,
    849622500, 849623400, 849624300, 849625200, 849626100, 849627000,
    849627900, 849628800, 849629700, 849630600, 849631500, 849632400,
    849633300, 849634200, 849635100, 849636000, 849636900, 849637800,
    849638700, 849639600, 849640500, 849641400, 849642300, 849643200,
    849644100, 849645000, 849645900, 849646800, 849647700, 849648600,
    849649500, 849650400, 849651300, 849652200, 849653100, 849654000,
    849654900, 849655800, 849656700, 849657600, 849658500, 849659400,
    849660300, 849661200, 849662100, 849663000, 849663900, 849664800,
    849665700, 849666600, 849667500, 849668400, 849669300, 849670200,
    849671100, 849672000, 849672900, 849673800, 849674700, 849675600,
    849676500, 849677400, 849678300, 849679200, 849680100, 849681000,
    849681900, 849682800, 849683700, 849684600, 849685500, 849686400,
    849687300, 849688200, 849689100, 849690000, 849690900, 849691800,
    849692700, 849693600, 849694500, 849695400, 849696300, 849697200,
    849698100, 849699000, 849699900, 849700800, 849701700, 849702600,
    849703500, 849704400, 849705300, 849706200, 849707100, 849708000,
    849708900, 849709800, 849710700, 849711600, 849712500, 849713400,
    849714300, 849715200, 849716100, 849717000, 849717900, 849718800,
    849719700, 849720600, 849721500, 849722400, 849723300, 849724200,
    849725100, 849726000, 849726900, 849727800, 849728700, 849729600,
    849730500, 849731400, 849732300, 849733200, 849734100, 849735000,
    849735900, 849736800, 849737700, 849738600, 849739500, 849740400,
    849741300, 849742200, 849743100, 849744000, 849744900, 849745800,
    849746700, 849747600, 849748500, 849749400, 849750300, 849751200,
    849752100, 849753000, 849753900, 849754800, 849755700, 849756600,
    849757500, 849758400, 849759300, 849760200, 849761100, 849762000,
    849762900, 849763800, 849764700, 849765600, 849766500, 849767400,
    849768300, 849769200, 849770100, 849771000, 849771900, 849772800,
    849773700, 849774600, 849775500, 849776400, 849777300, 849778200,
    849779100, 849780000, 849780900, 849781800, 849782700, 849783600,
    849784500, 849785400, 849786300, 849787200, 849788100, 849789000,
    849789900, 849790800, 849791700, 849792600, 849793500, 849794400,
    849795300, 849796200, 849797100, 849798000, 849798900, 849799800,
    849800700, 849801600, 849802500, 849803400, 849804300, 849805200,
    849806100, 849807000, 849807900, 849808800, 849809700, 849810600,
    849811500, 849812400, 849813300, 849814200, 849815100, 849816000,
    849816900, 849817800, 849818700, 849819600, 849820500, 849821400,
    849822300, 849823200, 849824100, 849825000, 849825900, 849826800,
    849827700, 849828600, 849829500, 849830400, 849831300, 849832200,
    849833100, 849834000, 849834900, 849835800, 849836700, 849837600,
    849838500, 849839400, 849840300, 849841200, 849842100, 849843000,
    849843900, 849844800, 849845700, 849846600, 849847500, 849848400,
    849849300, 849850200, 849851100, 849852000, 849852900, 849853800,
    849854700, 849855600, 849856500, 849857400, 849858300, 849859200,
    849860100, 849861000, 849861900, 849862800, 849863700, 849864600,
    849865500, 849866400, 849867300, 849868200, 849869100, 849870000,
    849870900, 849871800, 849872700, 849873600, 849874500, 849875400,
    849876300, 849877200, 849878100, 849879000, 849879900, 849880800,
    849881700, 849882600, 849883500, 849884400, 849885300, 849886200,
    849887100, 849888000, 849888900, 849889800, 849890700, 849891600,
    849892500, 849893400, 849894300, 849895200, 849896100, 849897000,
    849897900, 849898800, 849899700, 849900600, 849901500, 849902400,
    849903300, 849904200, 849905100, 849906000, 849906900, 849907800,
    849908700, 849909600, 849910500, 849911400, 849912300, 849913200,
    849914100, 849915000, 849915900, 849916800, 849917700, 849918600,
    849919500, 849920400, 849921300, 849922200, 849923100, 849924000,
    849924900, 849925800, 849926700, 849927600, 849928500, 849929400,
    849930300, 849931200, 849932100, 849933000, 849933900, 849934800,
    849935700, 849936600, 849937500, 849938400, 849939300, 849940200,
    849941100, 849942000, 849942900, 849943800, 849944700, 849945600,
    849946500, 849947400, 849948300, 849949200, 849950100, 849951000,
    849951900, 849952800, 849953700, 849954600, 849955500, 849956400,
    849957300, 849958200, 849959100, 849960000, 849960900, 849961800,
    849962700, 849963600, 849964500, 849965400, 849966300, 849967200,
    849968100, 849969000, 849969900, 849970800, 849971700, 849972600,
    849973500, 849974400, 849975300, 849976200, 849977100, 849978000,
    849978900, 849979800, 849980700, 849981600, 849982500, 849983400,
    849984300, 849985200, 849986100, 849987000, 849987900, 849988800,
    849989700, 849990600, 849991500, 849992400, 849993300, 849994200,
    849995100, 849996000, 849996900, 849997800, 849998700, 849999600,
    850000500, 850001400, 850002300, 850003200, 850004100, 850005000,
    850005900, 850006800, 850007700, 850008600, 850009500, 850010400,
    850011300, 850012200, 850013100, 850014000, 850014900, 850015800,
    850016700, 850017600, 850018500, 850019400, 850020300, 850021200,
    850022100, 850023000, 850023900, 850024800, 850025700, 850026600,
    850027500, 850028400, 850029300, 850030200, 850031100, 850032000,
    850032900, 850033800, 850034700, 850035600, 850036500, 850037400,
    850038300, 850039200, 850040100, 850041000, 850041900, 850042800,
    850043700, 850044600, 850045500, 850046400, 850047300, 850048200,
    850049100, 850050000, 850050900, 850051800, 850052700, 850053600,
    850054500, 850055400, 850056300, 850057200, 850058100, 850059000,
    850059900, 850060800, 850061700, 850062600, 850063500, 850064400,
    850065300, 850066200, 850067100, 850068000, 850068900, 850069800,
    850070700, 850071600, 850072500, 850073400, 850074300, 850075200,
    850076100, 850077000, 850077900, 850078800, 850079700, 850080600,
    850081500, 850082400, 850083300, 850084200, 850085100, 850086000,
    850086900, 850087800, 850088700, 850089600, 850090500, 850091400,
    850092300, 850093200, 850094100, 850095000, 850095900, 850096800,
    850097700, 850098600, 850099500, 850100400, 850101300, 850102200,
    850103100, 850104000, 850104900, 850105800, 850106700, 850107600,
    850108500, 850109400, 850110300, 850111200, 850112100, 850113000,
    850113900, 850114800, 850115700, 850116600, 850117500, 850118400,
    850119300, 850120200, 850121100, 850122000, 850122900, 850123800,
    850124700, 850125600, 850126500, 850127400, 850128300, 850129200,
    850130100, 850131000, 850131900, 850132800, 850133700, 850134600,
    850135500, 850136400, 850137300, 850138200, 850139100, 850140000,
    850140900, 850141800, 850142700, 850143600, 850144500, 850145400,
    850146300, 850147200, 850148100, 850149000, 850149900, 850150800,
    850151700, 850152600, 850153500, 850154400, 850155300, 850156200,
    850157100, 850158000, 850158900, 850159800, 850160700, 850161600,
    850162500, 850163400, 850164300, 850165200, 850166100, 850167000,
    850167900, 850168800, 850169700, 850170600, 850171500, 850172400,
    850173300, 850174200, 850175100, 850176000, 850176900, 850177800,
    850178700, 850179600, 850180500, 850181400, 850182300, 850183200,
    850184100, 850185000, 850185900, 850186800, 850187700, 850188600,
    850189500, 850190400, 850191300, 850192200, 850193100, 850194000,
    850194900, 850195800, 850196700, 850197600, 850198500, 850199400,
    850200300, 850201200, 850202100, 850203000, 850203900, 850204800,
    850205700, 850206600, 850207500, 850208400, 850209300, 850210200,
    850211100, 850212000, 850212900, 850213800, 850214700, 850215600,
    850216500, 850217400, 850218300, 850219200, 850220100, 850221000,
    850221900, 850222800, 850223700, 850224600, 850225500, 850226400,
    850227300, 850228200, 850229100, 850230000, 850230900, 850231800,
    850232700, 850233600, 850234500, 850235400, 850236300, 850237200,
    850238100, 850239000, 850239900, 850240800, 850241700, 850242600,
    850243500, 850244400, 850245300, 850246200, 850247100, 850248000,
    850248900, 850249800, 850250700, 850251600, 850252500, 850253400,
    850254300, 850255200, 850256100, 850257000, 850257900, 850258800,
    850259700, 850260600, 850261500, 850262400, 850263300, 850264200,
    850265100, 850266000, 850266900, 850267800, 850268700, 850269600,
    850270500, 850271400, 850272300, 850273200, 850274100, 850275000,
    850275900, 850276800, 850277700, 850278600, 850279500, 850280400,
    850281300, 850282200, 850283100, 850284000, 850284900, 850285800,
    850286700, 850287600, 850288500, 850289400, 850290300, 850291200,
    850292100, 850293000, 850293900, 850294800, 850295700, 850296600,
    850297500, 850298400, 850299300, 850300200, 850301100, 850302000,
    850302900, 850303800, 850304700, 850305600, 850306500, 850307400,
    850308300, 850309200, 850310100, 850311000, 850311900, 850312800,
    850313700, 850314600, 850315500, 850316400, 850317300, 850318200,
    850319100, 850320000, 850320900, 850321800, 850322700, 850323600,
    850324500, 850325400, 850326300, 850327200, 850328100, 850329000,
    850329900, 850330800, 850331700, 850332600, 850333500, 850334400,
    850335300, 850336200, 850337100, 850338000, 850338900, 850339800,
    850340700, 850341600, 850342500, 850343400, 850344300, 850345200,
    850346100, 850347000, 850347900, 850348800, 850349700, 850350600,
    850351500, 850352400, 850353300, 850354200, 850355100, 850356000,
    850356900, 850357800, 850358700, 850359600, 850360500, 850361400,
    850362300, 850363200, 850364100, 850365000, 850365900, 850366800,
    850367700, 850368600, 850369500, 850370400, 850371300, 850372200,
    850373100, 850374000, 850374900, 850375800, 850376700, 850377600,
    850378500, 850379400, 850380300, 850381200, 850382100, 850383000,
    850383900, 850384800, 850385700, 850386600, 850387500, 850388400,
    850389300, 850390200, 850391100, 850392000, 850392900, 850393800,
    850394700, 850395600, 850396500, 850397400, 850398300, 850399200,
    850400100, 850401000, 850401900, 850402800, 850403700, 850404600,
    850405500, 850406400, 850407300, 850408200, 850409100, 850410000,
    850410900, 850411800, 850412700, 850413600, 850414500, 850415400,
    850416300, 850417200, 850418100, 850419000, 850419900, 850420800,
    850421700, 850422600, 850423500, 850424400, 850425300, 850426200,
    850427100, 850428000, 850428900, 850429800, 850430700, 850431600,
    850432500, 850433400, 850434300, 850435200, 850436100, 850437000,
    850437900, 850438800, 850439700, 850440600, 850441500, 850442400,
    850443300, 850444200, 850445100, 850446000, 850446900, 850447800,
    850448700, 850449600, 850450500, 850451400, 850452300, 850453200,
    850454100, 850455000, 850455900, 850456800, 850457700, 850458600,
    850459500, 850460400, 850461300, 850462200, 850463100, 850464000,
    850464900, 850465800, 850466700, 850467600, 850468500, 850469400,
    850470300, 850471200, 850472100, 850473000, 850473900, 850474800,
    850475700, 850476600, 850477500, 850478400, 850479300, 850480200,
    850481100, 850482000, 850482900, 850483800, 850484700, 850485600,
    850486500, 850487400, 850488300, 850489200, 850490100, 850491000,
    850491900, 850492800, 850493700, 850494600, 850495500, 850496400,
    850497300, 850498200, 850499100, 850500000, 850500900, 850501800,
    850502700, 850503600, 850504500, 850505400, 850506300, 850507200,
    850508100, 850509000, 850509900, 850510800, 850511700, 850512600,
    850513500, 850514400, 850515300, 850516200, 850517100, 850518000,
    850518900, 850519800, 850520700, 850521600, 850522500, 850523400,
    850524300, 850525200, 850526100, 850527000, 850527900, 850528800,
    850529700, 850530600, 850531500, 850532400, 850533300, 850534200,
    850535100, 850536000, 850536900, 850537800, 850538700, 850539600,
    850540500, 850541400, 850542300, 850543200, 850544100, 850545000,
    850545900, 850546800, 850547700, 850548600, 850549500, 850550400,
    850551300, 850552200, 850553100, 850554000, 850554900, 850555800,
    850556700, 850557600, 850558500, 850559400, 850560300, 850561200,
    850562100, 850563000, 850563900, 850564800, 850565700, 850566600,
    850567500, 850568400, 850569300, 850570200, 850571100, 850572000,
    850572900, 850573800, 850574700, 850575600, 850576500, 850577400,
    850578300, 850579200, 850580100, 850581000, 850581900, 850582800,
    850583700, 850584600, 850585500, 850586400, 850587300, 850588200,
    850589100, 850590000, 850590900, 850591800, 850592700, 850593600,
    850616100, 850617000, 850617900, 850618800, 850619700, 850620600,
    850621500, 850622400, 850623300, 850624200, 850625100, 850626000,
    850626900, 850627800, 850628700, 850629600, 850630500, 850631400,
    850632300, 850633200, 850634100, 850635000, 850635900, 850636800,
    850637700, 850638600, 850639500, 850640400, 850641300, 850642200,
    850643100, 850644000, 850644900, 850645800, 850646700, 850647600,
    850648500, 850649400, 850650300, 850651200, 850652100, 850653000,
    850653900, 850654800, 850655700, 850656600, 850657500, 850658400,
    850659300, 850660200, 850661100, 850662000, 850662900, 850663800,
    850664700, 850665600, 850666500, 850667400, 850668300, 850669200,
    850670100, 850671000, 850671900, 850672800, 850673700, 850674600,
    850675500, 850676400, 850677300, 850678200, 850679100, 850680000,
    850680900, 850681800, 850682700, 850683600, 850684500, 850685400,
    850686300, 850687200, 850688100, 850689000, 850689900, 850690800,
    850691700, 850692600, 850693500, 850694400, 850695300, 850696200,
    850697100, 850698000, 850698900, 850699800, 850700700, 850701600,
    850702500, 850703400, 850704300, 850705200, 850706100, 850707000,
    850707900, 850708800, 850709700, 850710600, 850711500, 850712400,
    850713300, 850714200, 850715100, 850716000, 850716900, 850717800,
    850718700, 850719600, 850720500, 850721400, 850722300, 850723200,
    850724100, 850725000, 850725900, 850726800, 850727700, 850728600,
    850729500, 850730400, 850731300, 850732200, 850733100, 850734000,
    850734900, 850735800, 850736700, 850737600, 850738500, 850739400,
    850740300, 850741200, 850742100, 850743000, 850743900, 850744800,
    850745700, 850746600, 850747500, 850748400, 850749300, 850750200,
    850751100, 850752000, 850752900, 850753800, 850754700, 850755600,
    850756500, 850757400, 850758300, 850759200, 850760100, 850761000,
    850761900, 850762800, 850763700, 850764600, 850765500, 850766400,
    850767300, 850768200, 850769100, 850770000, 850770900, 850771800,
    850772700, 850773600, 850774500, 850775400, 850776300, 850777200,
    850778100, 850779000, 850779900, 850780800, 850781700, 850782600,
    850783500, 850784400, 850785300, 850786200, 850787100, 850788000,
    850788900, 850789800, 850790700, 850791600, 850792500, 850793400,
    850794300, 850795200, 850796100, 850797000, 850797900, 850798800,
    850799700, 850800600, 850801500, 850802400, 850803300, 850804200,
    850805100, 850806000, 850806900, 850807800, 850808700, 850809600,
    850810500, 850811400, 850812300, 850813200, 850814100, 850815000,
    850815900, 850816800, 850817700, 850818600, 850819500, 850820400,
    850821300, 850822200, 850823100, 850824000, 850824900, 850825800,
    850826700, 850827600, 850828500, 850829400, 850830300, 850831200,
    850832100, 850833000, 850833900, 850834800, 850835700, 850836600,
    850837500, 850838400, 850839300, 850840200, 850841100, 850842000,
    850842900, 850843800, 850844700, 850845600, 850846500, 850847400,
    850848300, 850849200, 850850100, 850851000, 850851900, 850852800,
    850853700, 850854600, 850855500, 850856400, 850857300, 850858200,
    850859100, 850860000, 850860900, 850861800, 850862700, 850863600,
    850864500, 850865400, 850866300, 850867200, 850868100, 850869000,
    850869900, 850870800, 850871700, 850872600, 850873500, 850874400,
    850875300, 850876200, 850877100, 850878000, 850878900, 850879800,
    850880700, 850881600, 850882500, 850883400, 850884300, 850885200,
    850886100, 850887000, 850887900, 850888800, 850889700, 850890600,
    850891500, 850892400, 850893300, 850894200, 850895100, 850896000,
    850896900, 850897800, 850898700, 850899600, 850900500, 850901400,
    850902300, 850903200, 850904100, 850905000, 850905900, 850906800,
    850907700, 850908600, 850909500, 850910400, 850911300, 850912200,
    850913100, 850914000, 850914900, 850915800, 850916700, 850917600,
    850918500, 850919400, 850920300, 850921200, 850922100, 850923000,
    850923900, 850924800, 850925700, 850926600, 850927500, 850928400,
    850929300, 850930200, 850931100, 850932000, 850932900, 850933800,
    850934700, 850935600, 850936500, 850937400, 850938300, 850939200,
    850940100, 850941000, 850941900, 850942800, 850943700, 850944600,
    850945500, 850946400, 850947300, 850948200, 850949100, 850950000,
    850950900, 850951800, 850952700, 850953600, 850954500, 850955400,
    850956300, 850957200, 850958100, 850959000, 850959900, 850960800,
    850961700, 850962600, 850963500, 850964400, 850965300, 850966200,
    850967100, 850968000, 850968900, 850969800, 850970700, 850971600,
    850972500, 850973400, 850974300, 850975200, 850976100, 850977000,
    850977900, 850978800, 850979700, 850980600, 850981500, 850982400,
    850983300, 850984200, 850985100, 850986000, 850986900, 850987800,
    850988700, 850989600, 850990500, 850991400, 850992300, 850993200,
    850994100, 850995000, 850995900, 850996800, 850997700, 850998600,
    850999500, 851000400, 851001300, 851002200, 851003100, 851004000,
    851004900, 851005800, 851006700, 851007600, 851008500, 851009400,
    851010300, 851011200, 851012100, 851013000, 851013900, 851014800,
    851015700, 851016600, 851017500, 851018400, 851019300, 851020200,
    851021100, 851022000, 851022900, 851023800, 851024700, 851025600,
    851026500, 851027400, 851028300, 851029200, 851030100, 851031000,
    851031900, 851032800, 851033700, 851034600, 851035500, 851036400,
    851037300, 851038200, 851039100, 851040000, 851040900, 851041800,
    851042700, 851043600, 851044500, 851045400, 851046300, 851047200,
    851048100, 851049000, 851049900, 851050800, 851051700, 851052600,
    851053500, 851054400, 851055300, 851056200, 851057100, 851058000,
    851058900, 851059800, 851060700, 851061600, 851062500, 851063400,
    851064300, 851065200, 851066100, 851067000, 851067900, 851068800,
    851069700, 851070600, 851071500, 851072400, 851073300, 851074200,
    851075100, 851076000, 851076900, 851077800, 851078700, 851079600,
    851080500, 851081400, 851082300, 851083200, 851084100, 851085000,
    851085900, 851086800, 851087700, 851088600, 851089500, 851090400,
    851091300, 851092200, 851093100, 851094000, 851094900, 851095800,
    851096700, 851097600, 851098500, 851099400, 851100300, 851101200,
    851102100, 851103000, 851103900, 851104800, 851105700, 851106600,
    851107500, 851108400, 851109300, 851110200, 851111100, 851112000,
    851112900, 851113800, 851114700, 851115600, 851116500, 851117400,
    851118300, 851119200, 851120100, 851121000, 851121900, 851122800,
    851123700, 851124600, 851125500, 851126400, 851127300, 851128200,
    851129100, 851130000, 851130900, 851131800, 851132700, 851133600,
    851134500, 851135400, 851136300, 851137200, 851138100, 851139000,
    851139900, 851140800, 851141700, 851142600, 851143500, 851144400,
    851145300, 851146200, 851147100, 851148000, 851148900, 851149800,
    851150700, 851151600, 851152500, 851153400, 851154300, 851155200,
    851156100, 851157000, 851157900, 851158800, 851159700, 851160600,
    851161500, 851162400, 851163300, 851164200, 851165100, 851166000,
    851166900, 851167800, 851168700, 851169600, 851170500, 851171400,
    851172300, 851173200, 851174100, 851175000, 851175900, 851176800,
    851177700, 851178600, 851179500, 851180400, 851181300, 851182200,
    851183100, 851184000, 851184900, 851185800, 851186700, 851187600,
    851188500, 851189400, 851190300, 851191200, 851192100, 851193000,
    851193900, 851194800, 851195700, 851196600, 851197500, 851198400,
    851199300, 851200200, 851201100, 851202000, 851202900, 851203800,
    851204700, 851205600, 851206500, 851207400, 851208300, 851209200,
    851210100, 851211000, 851211900, 851212800, 851213700, 851214600,
    851215500, 851216400, 851217300, 851218200, 851219100, 851220000,
    851220900, 851221800, 851222700, 851223600, 851224500, 851225400,
    851226300, 851227200, 851228100, 851229000, 851229900, 851230800,
    851231700, 851232600, 851233500, 851234400, 851235300, 851236200,
    851237100, 851238000, 851238900, 851239800, 851240700, 851241600,
    851242500, 851243400, 851244300, 851245200, 851246100, 851247000,
    851247900, 851248800, 851249700, 851250600, 851251500, 851252400,
    851253300, 851254200, 851255100, 851256000, 851256900, 851257800,
    851258700, 851259600, 851260500, 851261400, 851262300, 851263200,
    851264100, 851265000, 851265900, 851266800, 851267700, 851268600,
    851269500, 851270400, 851271300, 851272200, 851273100, 851274000,
    851274900, 851275800, 851276700, 851277600, 851278500, 851279400,
    851280300, 851281200, 851282100, 851283000, 851283900, 851284800,
    851285700, 851286600, 851287500, 851288400, 851289300, 851290200,
    851291100, 851292000, 851292900, 851293800, 851294700, 851295600,
    851296500, 851297400, 851298300, 851299200, 851300100, 851301000,
    851301900, 851302800, 851303700, 851304600, 851305500, 851306400,
    851307300, 851308200, 851309100, 851310000, 851310900, 851311800,
    851312700, 851313600, 851314500, 851315400, 851316300, 851317200,
    851318100, 851319000, 851319900, 851320800, 851321700, 851322600,
    851323500, 851324400, 851325300, 851326200, 851327100, 851328000,
    851328900, 851329800, 851330700, 851331600, 851332500, 851333400,
    851334300, 851335200, 851336100, 851337000, 851337900, 851338800,
    851339700, 851340600, 851341500, 851342400, 851343300, 851344200,
    851345100, 851346000, 851346900, 851347800, 851348700, 851349600,
    851350500, 851351400, 851352300, 851353200, 851354100, 851355000,
    851355900, 851356800, 851357700, 851358600, 851359500, 851360400,
    851361300, 851362200, 851363100, 851364000, 851364900, 851365800,
    851366700, 851367600, 851368500, 851369400, 851370300, 851371200,
    851372100, 851373000, 851373900, 851374800, 851375700, 851376600,
    851377500, 851378400, 851379300, 851380200, 851381100, 851382000,
    851382900, 851383800, 851384700, 851385600, 851386500, 851387400,
    851388300, 851389200, 851390100, 851391000, 851391900, 851392800,
    851393700, 851394600, 851395500, 851396400, 851397300, 851398200,
    851399100, 851400000, 851400900, 851401800, 851402700, 851403600,
    851404500, 851405400, 851406300, 851407200, 851408100, 851409000,
    851409900, 851410800, 851411700, 851412600, 851413500, 851414400,
    851415300, 851416200, 851417100, 851418000, 851418900, 851419800,
    851420700, 851421600, 851422500, 851423400, 851424300, 851425200,
    851426100, 851427000, 851427900, 851428800, 851429700, 851430600,
    851431500, 851432400, 851433300, 851434200, 851435100, 851436000,
    851436900, 851437800, 851438700, 851439600, 851440500, 851441400,
    851442300, 851443200, 851444100, 851445000, 851445900, 851446800,
    851447700, 851448600, 851449500, 851450400, 851451300, 851452200,
    851453100, 851454000, 851454900, 851455800, 851456700, 851457600,
    851458500, 851459400, 851460300, 851461200, 851462100, 851463000,
    851463900, 851464800, 851465700, 851466600, 851467500, 851468400,
    851469300, 851470200, 851471100, 851472000, 851472900, 851473800,
    851474700, 851475600, 851476500, 851477400, 851478300, 851479200,
    851480100, 851481000, 851481900, 851482800, 851483700, 851484600,
    851485500, 851486400, 851487300, 851488200, 851489100, 851490000,
    851490900, 851491800, 851492700, 851493600, 851494500, 851495400,
    851496300, 851497200, 851498100, 851499000, 851499900, 851500800,
    851501700, 851502600, 851503500, 851504400, 851505300, 851506200,
    851507100, 851508000, 851508900, 851509800, 851510700, 851511600,
    851512500, 851513400, 851514300, 851515200, 851516100, 851517000,
    851517900, 851518800, 851519700, 851520600, 851521500, 851522400,
    851523300, 851524200, 851525100, 851526000, 851526900, 851527800,
    851528700, 851529600, 851530500, 851531400, 851532300, 851533200,
    851534100, 851535000, 851535900, 851536800, 851537700, 851538600,
    851539500, 851540400, 851541300, 851542200, 851543100, 851544000,
    851544900, 851545800, 851546700, 851547600, 851548500, 851549400,
    851550300, 851551200, 851552100, 851553000, 851553900, 851554800,
    851555700, 851556600, 851557500, 851558400, 851559300, 851560200,
    851561100, 851562000, 851562900, 851563800, 851564700, 851565600,
    851566500, 851567400, 851568300, 851569200, 851570100, 851571000,
    851571900, 851572800, 851573700, 851574600, 851575500, 851576400,
    851577300, 851578200, 851579100, 851580000, 851580900, 851581800,
    851582700, 851583600, 851584500, 851585400, 851586300, 851587200,
    851588100, 851589000, 851589900, 851590800, 851591700, 851592600,
    851593500, 851594400, 851595300, 851596200, 851597100, 851598000,
    851598900, 851599800, 851600700, 851601600, 851602500, 851603400,
    851604300, 851605200, 851606100, 851607000, 851607900, 851608800,
    851609700, 851610600, 851611500, 851612400, 851613300, 851614200,
    851615100, 851616000, 851616900, 851617800, 851618700, 851619600,
    851620500, 851621400, 851622300, 851623200, 851624100, 851625000,
    851625900, 851626800, 851627700, 851628600, 851629500, 851630400,
    851631300, 851632200, 851633100, 851634000, 851634900, 851635800,
    851636700, 851637600, 851638500, 851639400, 851640300, 851641200,
    851642100, 851643000, 851643900, 851644800, 851645700, 851646600,
    851647500, 851648400, 851649300, 851650200, 851651100, 851652000,
    851652900, 851653800, 851654700, 851655600, 851656500, 851657400,
    851658300, 851659200, 851660100, 851661000, 851661900, 851662800,
    851663700, 851664600, 851665500, 851666400, 851667300, 851668200,
    851669100, 851670000, 851670900, 851671800, 851672700, 851673600,
    851674500, 851675400, 851676300, 851677200, 851678100, 851679000,
    851679900, 851680800, 851681700, 851682600, 851683500, 851684400,
    851685300, 851686200, 851687100, 851688000, 851688900, 851689800,
    851690700, 851691600, 851692500, 851693400, 851694300, 851695200,
    851696100, 851697000, 851697900, 851698800, 851699700, 851700600,
    851701500, 851702400, 851703300, 851704200, 851705100, 851706000,
    851706900, 851707800, 851708700, 851709600, 851710500, 851711400,
    851712300, 851713200, 851714100, 851715000, 851715900, 851716800,
    851717700, 851718600, 851719500, 851720400, 851721300, 851722200,
    851723100, 851724000, 851724900, 851725800, 851726700, 851727600,
    851728500, 851729400, 851730300, 851731200, 851732100, 851733000,
    851733900, 851734800, 851735700, 851736600, 851737500, 851738400,
    851739300, 851740200, 851741100, 851742000, 851742900, 851743800,
    851744700, 851745600, 851746500, 851747400, 851748300, 851749200,
    851750100, 851751000, 851751900, 851752800, 851753700, 851754600,
    851755500, 851756400, 851757300, 851758200, 851759100, 851760000,
    851760900, 851761800, 851762700, 851763600, 851764500, 851765400,
    851766300, 851767200, 851768100, 851769000, 851769900, 851770800,
    851771700, 851772600, 851773500, 851774400, 851775300, 851776200,
    851777100, 851778000, 851778900, 851779800, 851780700, 851781600,
    851782500, 851783400, 851784300, 851785200, 851786100, 851787000,
    851787900, 851788800, 851789700, 851790600, 851791500, 851792400,
    851793300, 851794200, 851795100, 851796000, 851796900, 851797800,
    851798700, 851799600, 851800500, 851801400, 851802300, 851803200,
    851804100, 851805000, 851805900, 851806800, 851807700, 851808600,
    851809500, 851810400, 851811300, 851812200, 851813100, 851814000,
    851814900, 851815800, 851816700, 851817600, 851818500, 851819400,
    851820300, 851821200, 851822100, 851823000, 851823900, 851824800,
    851825700, 851826600, 851827500, 851828400, 851829300, 851830200,
    851831100, 851832000, 851832900, 851833800, 851834700, 851835600,
    851836500, 851837400, 851838300, 851839200, 851840100, 851841000,
    851841900, 851842800, 851843700, 851844600, 851845500, 851846400,
    851847300, 851848200, 851849100, 851850000, 851850900, 851851800,
    851852700, 851853600, 851854500, 851855400, 851856300, 851857200,
    851858100, 851859000, 851859900, 851860800, 851861700, 851862600,
    851863500, 851864400, 851865300, 851866200, 851867100, 851868000,
    851868900, 851869800, 851870700, 851871600, 851872500, 851873400,
    851874300, 851875200, 851876100, 851877000, 851877900, 851878800,
    851879700, 851880600, 851881500, 851882400, 851883300, 851884200,
    851885100, 851886000, 851886900, 851887800, 851888700, 851889600,
    851890500, 851891400, 851892300, 851893200, 851894100, 851895000,
    851895900, 851896800, 851897700, 851898600, 851899500, 851900400,
    851901300, 851902200, 851903100, 851904000, 851904900, 851905800,
    851906700, 851907600, 851908500, 851909400, 851910300, 851911200,
    851912100, 851913000, 851913900, 851914800, 851915700, 851916600,
    851917500, 851918400, 851919300, 851920200, 851921100, 851922000,
    851922900, 851923800, 851924700, 851925600, 851926500, 851927400,
    851928300, 851929200, 851930100, 851931000, 851931900, 851932800,
    851933700, 851934600, 851935500, 851936400, 851937300, 851938200,
    851939100, 851940000, 851940900, 851941800, 851942700, 851943600,
    851944500, 851945400, 851946300, 851947200, 851948100, 851949000,
    851949900, 851950800, 851951700, 851952600, 851953500, 851954400,
    851955300, 851956200, 851957100, 851958000, 851958900, 851959800,
    851960700, 851961600, 851962500, 851963400, 851964300, 851965200,
    851966100, 851967000, 851967900, 851968800, 851969700, 851970600,
    851971500, 851972400, 851973300, 851974200, 851975100, 851976000,
    851976900, 851977800, 851978700, 851979600, 851980500, 851981400,
    851982300, 851983200, 851984100, 851985000, 851985900, 851986800,
    851987700, 851988600, 851989500, 851990400, 851991300, 851992200,
    851993100, 851994000, 851994900, 851995800, 851996700, 851997600,
    851998500, 851999400, 852000300, 852001200, 852002100, 852003000,
    852003900, 852004800, 852005700, 852006600, 852007500, 852008400,
    852009300, 852010200, 852011100, 852012000, 852012900, 852013800,
    852014700, 852015600, 852016500, 852017400, 852018300, 852019200,
    852020100, 852021000, 852021900, 852022800, 852023700, 852024600,
    852025500, 852026400, 852027300, 852028200, 852029100, 852030000,
    852030900, 852031800, 852032700, 852033600, 852034500, 852035400,
    852036300, 852037200, 852038100, 852039000, 852039900, 852040800,
    852041700, 852042600, 852043500, 852044400, 852045300, 852046200,
    852047100, 852048000, 852048900, 852049800, 852050700, 852051600,
    852052500, 852053400, 852054300, 852055200, 852056100, 852057000,
    852057900, 852058800, 852059700, 852060600, 852061500, 852062400,
    852063300, 852064200, 852065100, 852066000, 852066900, 852067800,
    852068700, 852069600, 852070500, 852071400, 852072300, 852073200,
    852074100, 852075000, 852075900, 852076800, 852077700, 852078600,
    852079500, 852080400, 852081300, 852082200, 852083100, 852084000,
    852084900, 852085800, 852086700, 852087600, 852088500, 852089400,
    852090300, 852091200, 852092100, 852093000, 852093900, 852094800,
    852095700, 852096600, 852097500, 852098400, 852099300, 852100200,
    852101100, 852102000, 852102900, 852103800, 852104700, 852105600,
    852106500, 852107400, 852108300, 852109200, 852110100, 852111000,
    852111900, 852112800, 852113700, 852114600, 852115500, 852116400,
    852117300, 852118200, 852119100, 852120000, 852120900, 852121800,
    852122700, 852123600, 852124500, 852125400, 852126300, 852127200,
    852128100, 852129000, 852129900, 852130800, 852131700, 852132600,
    852133500, 852134400, 852135300, 852136200, 852137100, 852138000,
    852138900, 852139800, 852140700, 852141600, 852142500, 852143400,
    852144300, 852145200, 852146100, 852147000, 852147900, 852148800,
    852149700, 852150600, 852151500, 852152400, 852153300, 852154200,
    852155100, 852156000, 852156900, 852157800, 852158700, 852159600,
    852160500, 852161400, 852162300, 852163200, 852164100, 852165000,
    852165900, 852166800, 852167700, 852168600, 852169500, 852170400,
    852171300, 852172200, 852173100, 852174000, 852174900, 852175800,
    852176700, 852177600, 852178500, 852179400, 852180300, 852181200,
    852182100, 852183000, 852183900, 852184800, 852185700, 852186600,
    852187500, 852188400, 852189300, 852190200, 852191100, 852192000,
    852192900, 852193800, 852194700, 852195600, 852196500, 852197400,
    852198300, 852199200, 852200100, 852201000, 852201900, 852202800,
    852203700, 852204600, 852205500, 852206400, 852207300, 852208200,
    852209100, 852210000, 852210900, 852211800, 852212700, 852213600,
    852214500, 852215400, 852216300, 852217200, 852218100, 852219000,
    852219900, 852220800, 852221700, 852222600, 852223500, 852224400,
    852225300, 852226200, 852227100, 852228000, 852228900, 852229800,
    852230700, 852231600, 852232500, 852233400, 852234300, 852235200,
    852236100, 852237000, 852237900, 852238800, 852239700, 852240600,
    852241500, 852242400, 852243300, 852244200, 852245100, 852246000,
    852246900, 852247800, 852248700, 852249600, 852250500, 852251400,
    852252300, 852253200, 852254100, 852255000, 852255900, 852256800,
    852257700, 852258600, 852259500, 852260400, 852261300, 852262200,
    852263100, 852264000, 852264900, 852265800, 852266700, 852267600,
    852268500, 852269400, 852270300, 852271200, 852272100, 852273000,
    852273900, 852274800, 852275700, 852276600, 852277500, 852278400,
    852279300, 852280200, 852281100, 852282000, 852282900, 852283800,
    852284700, 852285600, 852286500, 852287400, 852288300, 852289200,
    852290100, 852291000, 852291900, 852292800, 852293700, 852294600,
    852295500, 852296400, 852297300, 852298200, 852299100, 852300000,
    852300900, 852301800, 852302700, 852303600, 852304500, 852305400,
    852306300, 852307200, 852308100, 852309000, 852309900, 852310800,
    852311700, 852312600, 852313500, 852314400, 852315300, 852316200,
    852317100, 852318000, 852318900, 852319800, 852320700, 852321600,
    852322500, 852323400, 852324300, 852325200, 852326100, 852327000,
    852327900, 852328800, 852329700, 852330600, 852331500, 852332400,
    852333300, 852334200, 852335100, 852336000, 852336900, 852337800,
    852338700, 852339600, 852340500, 852341400, 852342300, 852343200,
    852344100, 852345000, 852345900, 852346800, 852347700, 852348600,
    852349500, 852350400, 852351300, 852352200, 852353100, 852354000,
    852354900, 852355800, 852356700, 852357600, 852358500, 852359400,
    852360300, 852361200, 852362100, 852363000, 852363900, 852364800,
    852365700, 852366600, 852367500, 852368400, 852369300, 852370200,
    852371100, 852372000, 852372900, 852373800, 852374700, 852375600,
    852376500, 852377400, 852378300, 852379200, 852380100, 852381000,
    852381900, 852382800, 852383700, 852384600, 852385500, 852386400,
    852387300, 852388200, 852389100, 852390000, 852390900, 852391800,
    852392700, 852393600, 852394500, 852395400, 852396300, 852397200,
    852398100, 852399000, 852399900, 852400800, 852401700, 852402600,
    852403500, 852404400, 852405300, 852406200, 852407100, 852408000,
    852408900, 852409800, 852410700, 852411600, 852412500, 852413400,
    852414300, 852415200, 852416100, 852417000, 852417900, 852418800,
    852419700, 852420600, 852421500, 852422400, 852423300, 852424200,
    852425100, 852426000, 852426900, 852427800, 852428700, 852429600,
    852430500, 852431400, 852432300, 852433200, 852434100, 852435000,
    852435900, 852436800, 852437700, 852438600, 852439500, 852440400,
    852441300, 852442200, 852443100, 852444000, 852444900, 852445800,
    852446700, 852447600, 852448500, 852449400, 852450300, 852451200,
    852452100, 852453000, 852453900, 852454800, 852455700, 852456600,
    852457500, 852458400, 852459300, 852460200, 852461100, 852462000,
    852462900, 852463800, 852464700, 852465600, 852466500, 852467400,
    852468300, 852469200, 852470100, 852471000, 852471900, 852472800,
    852473700, 852474600, 852475500, 852476400, 852477300, 852478200,
    852479100, 852480000, 852480900, 852481800, 852482700, 852483600,
    852484500, 852485400, 852486300, 852487200, 852488100, 852489000,
    852489900, 852490800, 852491700, 852492600, 852493500, 852494400,
    852495300, 852496200, 852497100, 852498000, 852498900, 852499800,
    852500700, 852501600, 852502500, 852503400, 852504300, 852505200,
    852506100, 852507000, 852507900, 852508800, 852509700, 852510600,
    852511500, 852512400, 852513300, 852514200, 852515100, 852516000,
    852516900, 852517800, 852518700, 852519600, 852520500, 852521400,
    852522300, 852523200, 852524100, 852525000, 852525900, 852526800,
    852527700, 852528600, 852529500, 852530400, 852531300, 852532200,
    852533100, 852534000, 852534900, 852535800, 852536700, 852537600,
    852538500, 852539400, 852540300, 852541200, 852542100, 852543000,
    852543900, 852544800, 852545700, 852546600, 852547500, 852548400,
    852549300, 852550200, 852551100, 852552000, 852552900, 852553800,
    852554700, 852555600, 852556500, 852557400, 852558300, 852559200,
    852560100, 852561000, 852561900, 852562800, 852563700, 852564600,
    852565500, 852566400, 852567300, 852568200, 852569100, 852570000,
    852570900, 852571800, 852572700, 852573600, 852574500, 852575400,
    852576300, 852577200, 852578100, 852579000, 852579900, 852580800,
    852581700, 852582600, 852583500, 852584400, 852585300, 852586200,
    852587100, 852588000, 852588900, 852589800, 852590700, 852591600,
    852592500, 852593400, 852594300, 852595200, 852596100, 852597000,
    852597900, 852598800, 852599700, 852600600, 852601500, 852602400,
    852603300, 852604200, 852605100, 852606000, 852606900, 852607800,
    852608700, 852609600, 852610500, 852611400, 852612300, 852613200,
    852614100, 852615000, 852615900, 852616800, 852617700, 852618600,
    852619500, 852620400, 852621300, 852622200, 852623100, 852624000,
    852624900, 852625800, 852626700, 852627600, 852628500, 852629400,
    852630300, 852631200, 852632100, 852633000, 852633900, 852634800,
    852635700, 852636600, 852637500, 852638400, 852639300, 852640200,
    852641100, 852642000, 852642900, 852643800, 852644700, 852645600,
    852646500, 852647400, 852648300, 852649200, 852650100, 852651000,
    852651900, 852652800, 852653700, 852654600, 852655500, 852656400,
    852657300, 852658200, 852659100, 852660000, 852660900, 852661800,
    852662700, 852663600, 852664500, 852665400, 852666300, 852667200,
    852668100, 852669000, 852669900, 852670800, 852671700, 852672600,
    852673500, 852674400, 852675300, 852676200, 852677100, 852678000,
    852678900, 852679800, 852680700, 852681600, 852682500, 852683400,
    852684300, 852685200, 852686100, 852687000, 852687900, 852688800,
    852689700, 852690600, 852691500, 852692400, 852693300, 852694200,
    852695100, 852696000, 852696900, 852697800, 852698700, 852699600,
    852700500, 852701400, 852702300, 852703200, 852704100, 852705000,
    852705900, 852706800, 852707700, 852708600, 852709500, 852710400,
    852711300, 852712200, 852713100, 852714000, 852714900, 852715800,
    852716700, 852717600, 852718500, 852719400, 852720300, 852721200,
    852722100, 852723000, 852723900, 852724800, 852725700, 852726600,
    852727500, 852728400, 852729300, 852730200, 852731100, 852732000,
    852732900, 852733800, 852734700, 852735600, 852736500, 852737400,
    852738300, 852739200, 852740100, 852741000, 852741900, 852742800,
    852743700, 852744600, 852745500, 852746400, 852747300, 852748200,
    852749100, 852750000, 852750900, 852751800, 852752700, 852753600,
    852754500, 852755400, 852756300, 852757200, 852758100, 852759000,
    852759900, 852760800, 852761700, 852762600, 852763500, 852764400,
    852765300, 852766200, 852767100, 852768000, 852768900, 852769800,
    852770700, 852771600, 852772500, 852773400, 852774300, 852775200,
    852776100, 852777000, 852777900, 852778800, 852779700, 852780600,
    852781500, 852782400, 852783300, 852784200, 852785100, 852786000,
    852786900, 852787800, 852788700, 852789600, 852790500, 852791400,
    852792300, 852793200, 852794100, 852795000, 852795900, 852796800,
    852797700, 852798600, 852799500, 852800400, 852801300, 852802200,
    852803100, 852804000, 852804900, 852805800, 852806700, 852807600,
    852808500, 852809400, 852810300, 852811200, 852812100, 852813000,
    852813900, 852814800, 852815700, 852816600, 852817500, 852818400,
    852819300, 852820200, 852821100, 852822000, 852822900, 852823800,
    852824700, 852825600, 852826500, 852827400, 852828300, 852829200,
    852830100, 852831000, 852831900, 852832800, 852833700, 852834600,
    852835500, 852836400, 852837300, 852838200, 852839100, 852840000,
    852840900, 852841800, 852842700, 852843600, 852844500, 852845400,
    852846300, 852847200, 852848100, 852849000, 852849900, 852850800,
    852851700, 852852600, 852853500, 852854400, 852855300, 852856200,
    852857100, 852858000, 852858900, 852859800, 852860700, 852861600,
    852862500, 852863400, 852864300, 852865200, 852866100, 852867000,
    852867900, 852868800, 852869700, 852870600, 852871500, 852872400,
    852873300, 852874200, 852875100, 852876000, 852876900, 852877800,
    852878700, 852879600, 852880500, 852881400, 852882300, 852883200,
    852884100, 852885000, 852885900, 852886800, 852887700, 852888600,
    852889500, 852890400, 852891300, 852892200, 852893100, 852894000,
    852894900, 852895800, 852896700, 852897600, 852898500, 852899400,
    852900300, 852901200, 852902100, 852903000, 852903900, 852904800,
    852905700, 852906600, 852907500, 852908400, 852909300, 852910200,
    852911100, 852912000, 852912900, 852913800, 852914700, 852915600,
    852916500, 852917400, 852918300, 852919200, 852920100, 852921000,
    852921900, 852922800, 852923700, 852924600, 852925500, 852926400,
    852927300, 852928200, 852929100, 852930000, 852930900, 852931800,
    852932700, 852933600, 852934500, 852935400, 852936300, 852937200,
    852938100, 852939000, 852939900, 852940800, 852941700, 852942600,
    852943500, 852944400, 852945300, 852946200, 852947100, 852948000,
    852948900, 852949800, 852950700, 852951600, 852952500, 852953400,
    852954300, 852955200, 852956100, 852957000, 852957900, 852958800,
    852959700, 852960600, 852961500, 852962400, 852963300, 852964200,
    852965100, 852966000, 852966900, 852967800, 852968700, 852969600,
    852970500, 852971400, 852972300, 852973200, 852974100, 852975000,
    852975900, 852976800, 852977700, 852978600, 852979500, 852980400,
    852981300, 852982200, 852983100, 852984000, 852984900, 852985800,
    852986700, 852987600, 852988500, 852989400, 852990300, 852991200,
    852992100, 852993000, 852993900, 852994800, 852995700, 852996600,
    852997500, 852998400, 852999300, 853000200, 853001100, 853002000,
    853002900, 853003800, 853004700, 853005600, 853006500, 853007400,
    853008300, 853009200, 853010100, 853011000, 853011900, 853012800,
    853013700, 853014600, 853015500, 853016400, 853017300, 853018200,
    853019100, 853020000, 853020900, 853021800, 853022700, 853023600,
    853024500, 853025400, 853026300, 853027200, 853028100, 853029000,
    853029900, 853030800, 853031700, 853032600, 853033500, 853034400,
    853035300, 853036200, 853037100, 853038000, 853038900, 853039800,
    853040700, 853041600, 853042500, 853043400, 853044300, 853045200,
    853046100, 853047000, 853047900, 853048800, 853049700, 853050600,
    853051500, 853052400, 853053300, 853054200, 853055100, 853056000,
    853056900, 853057800, 853058700, 853059600, 853060500, 853061400,
    853062300, 853063200, 853064100, 853065000, 853065900, 853066800,
    853067700, 853068600, 853069500, 853070400, 853071300, 853072200,
    853073100, 853074000, 853074900, 853075800, 853076700, 853077600,
    853078500, 853079400, 853080300, 853081200, 853082100, 853083000,
    853083900, 853084800, 853085700, 853086600, 853087500, 853088400,
    853089300, 853090200, 853091100, 853092000, 853092900, 853093800,
    853094700, 853095600, 853096500, 853097400, 853098300, 853099200,
    853100100, 853101000, 853101900, 853102800, 853103700, 853104600,
    853105500, 853106400, 853107300, 853108200, 853109100, 853110000,
    853110900, 853111800, 853112700, 853113600, 853114500, 853115400,
    853116300, 853117200, 853118100, 853119000, 853119900, 853120800,
    853121700, 853122600, 853123500, 853124400, 853125300, 853126200,
    853127100, 853128000, 853128900, 853129800, 853130700, 853131600,
    853132500, 853133400, 853134300, 853135200, 853136100, 853137000,
    853137900, 853138800, 853139700, 853140600, 853141500, 853142400,
    853143300, 853144200, 853145100, 853146000, 853146900, 853147800,
    853148700, 853149600, 853150500, 853151400, 853152300, 853153200,
    853154100, 853155000, 853155900, 853156800, 853157700, 853158600,
    853159500, 853160400, 853161300, 853162200, 853163100, 853164000,
    853164900, 853165800, 853166700, 853167600, 853168500, 853169400,
    853170300, 853171200, 853172100, 853173000, 853173900, 853174800,
    853175700, 853176600, 853177500, 853178400, 853179300, 853180200,
    853181100, 853182000, 853182900, 853183800, 853184700, 853185600,
    853186500, 853187400, 853188300, 853189200, 853190100, 853191000,
    853191900, 853192800, 853193700, 853194600, 853195500, 853196400,
    853197300, 853198200, 853199100, 853200000, 853200900, 853201800,
    853202700, 853203600, 853204500, 853205400, 853206300, 853207200,
    853208100, 853209000, 853209900, 853210800, 853211700, 853212600,
    853213500, 853214400, 853215300, 853216200, 853217100, 853218000,
    853218900, 853219800, 853220700, 853221600, 853222500, 853223400,
    853224300, 853225200, 853226100, 853227000, 853227900, 853228800,
    853229700, 853230600, 853231500, 853232400, 853233300, 853234200,
    853235100, 853236000, 853236900, 853237800, 853238700, 853239600,
    853240500, 853241400, 853242300, 853243200, 853244100, 853245000,
    853245900, 853246800, 853247700, 853248600, 853249500, 853250400,
    853251300, 853252200, 853253100, 853254000, 853254900, 853255800,
    853256700, 853257600, 853258500, 853259400, 853260300, 853261200,
    853262100, 853263000, 853263900, 853264800, 853265700, 853266600,
    853267500, 853268400, 853269300, 853270200, 853271100, 853272000,
    853272900, 853273800, 853274700, 853275600, 853276500, 853277400,
    853278300, 853279200, 853280100, 853281000, 853281900, 853282800,
    853283700, 853284600, 853285500, 853286400, 853287300, 853288200,
    853289100, 853290000, 853290900, 853291800, 853292700, 853293600,
    853294500, 853295400, 853296300, 853297200, 853298100, 853299000,
    853299900, 853300800, 853301700, 853302600, 853303500, 853304400,
    853305300, 853306200, 853307100, 853308000, 853308900, 853309800,
    853310700, 853311600, 853312500, 853313400, 853314300, 853315200,
    853316100, 853317000, 853317900, 853318800, 853319700, 853320600,
    853321500, 853322400, 853323300, 853324200, 853325100, 853326000,
    853326900, 853327800, 853328700, 853329600, 853330500, 853331400,
    853332300, 853333200, 853334100, 853335000, 853335900, 853336800,
    853337700, 853338600, 853339500, 853340400, 853341300, 853342200,
    853343100, 853344000, 853344900, 853345800, 853346700, 853347600,
    853348500, 853349400, 853350300, 853351200, 853352100, 853353000,
    853353900, 853354800, 853355700, 853356600, 853357500, 853358400,
    853359300, 853360200, 853361100, 853362000, 853362900, 853363800,
    853364700, 853365600, 853366500, 853367400, 853368300, 853369200,
    853370100, 853371000, 853371900, 853372800, 853373700, 853374600,
    853375500, 853376400, 853377300, 853378200, 853379100, 853380000,
    853380900, 853381800, 853382700, 853383600, 853384500, 853385400,
    853386300, 853387200, 853388100, 853389000, 853389900, 853390800,
    853391700, 853392600, 853393500, 853394400, 853395300, 853396200,
    853397100, 853398000, 853398900, 853399800, 853400700, 853401600,
    853402500, 853403400, 853404300, 853405200, 853406100, 853407000,
    853407900, 853408800, 853409700, 853410600, 853411500, 853412400,
    853413300, 853414200, 853415100, 853416000, 853416900, 853417800,
    853418700, 853419600, 853420500, 853421400, 853422300, 853423200,
    853424100, 853425000, 853425900, 853426800, 853427700, 853428600,
    853429500, 853430400, 853431300, 853432200, 853433100, 853434000,
    853434900, 853435800, 853436700, 853437600, 853438500, 853439400,
    853440300, 853441200, 853442100, 853443000, 853443900, 853444800,
    853445700, 853446600, 853447500, 853448400, 853449300, 853450200,
    853451100, 853452000, 853452900, 853453800, 853454700, 853455600,
    853456500, 853457400, 853458300, 853459200, 853460100, 853461000,
    853461900, 853462800, 853463700, 853464600, 853465500, 853466400,
    853467300, 853468200, 853469100, 853470000, 853470900, 853471800,
    853472700, 853473600, 853474500, 853475400, 853476300, 853477200,
    853478100, 853479000, 853479900, 853480800, 853481700, 853482600,
    853483500, 853484400, 853485300, 853486200, 853487100, 853488000,
    853488900, 853489800, 853490700, 853491600, 853492500, 853493400,
    853494300, 853495200, 853496100, 853497000, 853497900, 853498800,
    853499700, 853500600, 853501500, 853502400, 853503300, 853504200,
    853505100, 853506000, 853506900, 853507800, 853508700, 853509600,
    853510500, 853511400, 853512300, 853513200, 853514100, 853515000,
    853515900, 853516800, 853517700, 853518600, 853519500, 853520400,
    853521300, 853522200, 853523100, 853524000, 853524900, 853525800,
    853526700, 853527600, 853528500, 853529400, 853530300, 853531200,
    853532100, 853533000, 853533900, 853534800, 853535700, 853536600,
    853537500, 853538400, 853539300, 853540200, 853541100, 853542000,
    853542900, 853543800, 853544700, 853545600, 853546500, 853547400,
    853548300, 853549200, 853550100, 853551000, 853551900, 853552800,
    853553700, 853554600, 853555500, 853556400, 853557300, 853558200,
    853559100, 853560000, 853560900, 853561800, 853562700, 853563600,
    853564500, 853565400, 853566300, 853567200, 853568100, 853569000,
    853569900, 853570800, 853571700, 853572600, 853573500, 853574400,
    853575300, 853576200, 853577100, 853578000, 853578900, 853579800,
    853580700, 853581600, 853582500, 853583400, 853584300, 853585200,
    853586100, 853587000, 853587900, 853588800, 853589700, 853590600,
    853591500, 853592400, 853593300, 853594200, 853595100, 853596000,
    853596900, 853597800, 853598700, 853599600, 853600500, 853601400,
    853602300, 853603200, 853604100, 853605000, 853605900, 853606800,
    853607700, 853608600, 853609500, 853610400, 853611300, 853612200,
    853613100, 853614000, 853614900, 853615800, 853616700, 853617600,
    853618500, 853619400, 853620300, 853621200, 853622100, 853623000,
    853623900, 853624800, 853625700, 853626600, 853627500, 853628400,
    853629300, 853630200, 853631100, 853632000, 853632900, 853633800,
    853634700, 853635600, 853636500, 853637400, 853638300, 853639200,
    853640100, 853641000, 853641900, 853642800, 853643700, 853644600,
    853645500, 853646400, 853647300, 853648200, 853649100, 853650000,
    853650900, 853651800, 853652700, 853653600, 853654500, 853655400,
    853656300, 853657200, 853658100, 853659000, 853659900, 853660800,
    853661700, 853662600, 853663500, 853664400, 853665300, 853666200,
    853667100, 853668000, 853668900, 853669800, 853670700, 853671600,
    853672500, 853673400, 853674300, 853675200, 853676100, 853677000,
    853677900, 853678800, 853679700, 853680600, 853681500, 853682400,
    853683300, 853684200, 853685100, 853686000, 853686900, 853687800,
    853688700, 853689600, 853690500, 853691400, 853692300, 853693200,
    853694100, 853695000, 853695900, 853696800, 853697700, 853698600,
    853699500, 853700400, 853701300, 853702200, 853703100, 853704000,
    853704900, 853705800, 853706700, 853707600, 853708500, 853709400,
    853710300, 853711200, 853712100, 853713000, 853713900, 853714800,
    853715700, 853716600, 853717500, 853718400, 853719300, 853720200,
    853721100, 853722000, 853722900, 853723800, 853724700, 853725600,
    853726500, 853727400, 853728300, 853729200, 853730100, 853731000,
    853731900, 853732800, 853733700, 853734600, 853735500, 853736400,
    853737300, 853738200, 853739100, 853740000, 853740900, 853741800,
    853742700, 853743600, 853744500, 853745400, 853746300, 853747200,
    853748100, 853749000, 853749900, 853750800, 853751700, 853752600,
    853753500, 853754400, 853755300, 853756200, 853757100, 853758000,
    853758900, 853759800, 853760700, 853761600, 853762500, 853763400,
    853764300, 853765200, 853766100, 853767000, 853767900, 853768800,
    853769700, 853770600, 853771500, 853772400, 853773300, 853774200,
    853775100, 853776000, 853776900, 853777800, 853778700, 853779600,
    853780500, 853781400, 853782300, 853783200, 853784100, 853785000,
    853785900, 853786800, 853787700, 853788600, 853789500, 853790400,
    853791300, 853792200, 853793100, 853794000, 853794900, 853795800,
    853796700, 853797600, 853798500, 853799400, 853800300, 853801200,
    853802100, 853803000, 853803900, 853804800, 853805700, 853806600,
    853807500, 853808400, 853809300, 853810200, 853811100, 853812000,
    853812900, 853813800, 853814700, 853815600, 853816500, 853817400,
    853818300, 853819200, 853820100, 853821000, 853821900, 853822800,
    853823700, 853824600, 853825500, 853826400, 853827300, 853828200,
    853829100, 853830000, 853830900, 853831800, 853832700, 853833600,
    853834500, 853835400, 853836300, 853837200, 853838100, 853839000,
    853839900, 853840800, 853841700, 853842600, 853843500, 853844400,
    853845300, 853846200, 853847100, 853848000, 853848900, 853849800,
    853850700, 853851600, 853852500, 853853400, 853854300, 853855200,
    853856100, 853857000, 853857900, 853858800, 853859700, 853860600,
    853861500, 853862400, 853863300, 853864200, 853865100, 853866000,
    853866900, 853867800, 853868700, 853869600, 853870500, 853871400,
    853872300, 853873200, 853874100, 853875000, 853875900, 853876800,
    853877700, 853878600, 853879500, 853880400, 853881300, 853882200,
    853883100, 853884000, 853884900, 853885800, 853886700, 853887600,
    853888500, 853889400, 853890300, 853891200, 853892100, 853893000,
    853893900, 853894800, 853895700, 853896600, 853897500, 853898400,
    853899300, 853900200, 853901100, 853902000, 853902900, 853903800,
    853904700, 853905600, 853906500, 853907400, 853908300, 853909200,
    853910100, 853911000, 853911900, 853912800, 853913700, 853914600,
    853915500, 853916400, 853917300, 853918200, 853919100, 853920000,
    853920900, 853921800, 853922700, 853923600, 853924500, 853925400,
    853926300, 853927200, 853928100, 853929000, 853929900, 853930800,
    853931700, 853932600, 853933500, 853934400, 853935300, 853936200,
    853937100, 853938000, 853938900, 853939800, 853940700, 853941600,
    853942500, 853943400, 853944300, 853945200, 853946100, 853947000,
    853947900, 853948800, 853949700, 853950600, 853951500, 853952400,
    853953300, 853954200, 853955100, 853956000, 853956900, 853957800,
    853958700, 853959600, 853960500, 853961400, 853962300, 853963200,
    853964100, 853965000, 853965900, 853966800, 853967700, 853968600,
    853969500, 853970400, 853971300, 853972200, 853973100, 853974000,
    853974900, 853975800, 853976700, 853977600, 853978500, 853979400,
    853980300, 853981200, 853982100, 853983000, 853983900, 853984800,
    853985700, 853986600, 853987500, 853988400, 853989300, 853990200,
    853991100, 853992000, 853992900, 853993800, 853994700, 853995600,
    853996500, 853997400, 853998300, 853999200, 854000100, 854001000,
    854001900, 854002800, 854003700, 854004600, 854005500, 854006400,
    854007300, 854008200, 854009100, 854010000, 854010900, 854011800,
    854012700, 854013600, 854014500, 854015400, 854016300, 854017200,
    854018100, 854019000, 854019900, 854020800, 854021700, 854022600,
    854023500, 854024400, 854025300, 854026200, 854027100, 854028000,
    854028900, 854029800, 854030700, 854031600, 854032500, 854033400,
    854034300, 854035200, 854036100, 854037000, 854037900, 854038800,
    854039700, 854040600, 854041500, 854042400, 854043300, 854044200,
    854045100, 854046000, 854046900, 854047800, 854048700, 854049600,
    854050500, 854051400, 854052300, 854053200, 854054100, 854055000,
    854055900, 854056800, 854057700, 854058600, 854059500, 854060400,
    854061300, 854062200, 854063100, 854064000, 854064900, 854065800,
    854066700, 854067600, 854068500, 854069400, 854070300, 854071200,
    854072100, 854073000, 854073900, 854074800, 854075700, 854076600,
    854077500, 854078400, 854079300, 854080200, 854081100, 854082000,
    854082900, 854083800, 854084700, 854085600, 854086500, 854087400,
    854088300, 854089200, 854090100, 854091000, 854091900, 854092800,
    854093700, 854094600, 854095500, 854096400, 854097300, 854098200,
    854099100, 854100000, 854100900, 854101800, 854102700, 854103600,
    854104500, 854105400, 854106300, 854107200, 854108100, 854109000,
    854109900, 854110800, 854111700, 854112600, 854113500, 854114400,
    854115300, 854116200, 854117100, 854118000, 854118900, 854119800,
    854120700, 854121600, 854122500, 854123400, 854124300, 854125200,
    854126100, 854127000, 854127900, 854128800, 854129700, 854130600,
    854131500, 854132400, 854133300, 854134200, 854135100, 854136000,
    854136900, 854137800, 854138700, 854139600, 854140500, 854141400,
    854142300, 854143200, 854144100, 854145000, 854145900, 854146800,
    854147700, 854148600, 854149500, 854150400, 854151300, 854152200,
    854153100, 854154000, 854154900, 854155800, 854156700, 854157600,
    854158500, 854159400, 854160300, 854161200, 854162100, 854163000,
    854163900, 854164800, 854165700, 854166600, 854167500, 854168400,
    854169300, 854170200, 854171100, 854172000, 854172900, 854173800,
    854174700, 854175600, 854176500, 854177400, 854178300, 854179200,
    854180100, 854181000, 854181900, 854182800, 854183700, 854184600,
    854185500, 854186400, 854187300, 854188200, 854189100, 854190000,
    854190900, 854191800, 854192700, 854193600, 854194500, 854195400,
    854196300, 854197200, 854198100, 854199000, 854199900, 854200800,
    854201700, 854202600, 854203500, 854204400, 854205300, 854206200,
    854207100, 854208000, 854208900, 854209800, 854210700, 854211600,
    854212500, 854213400, 854214300, 854215200, 854216100, 854217000,
    854217900, 854218800, 854219700, 854220600, 854221500, 854222400,
    854223300, 854224200, 854225100, 854226000, 854226900, 854227800,
    854228700, 854229600, 854230500, 854231400, 854232300, 854233200,
    854234100, 854235000, 854235900, 854236800, 854237700, 854238600,
    854239500, 854240400, 854241300, 854242200, 854243100, 854244000,
    854244900, 854245800, 854246700, 854247600, 854248500, 854249400,
    854250300, 854251200, 854252100, 854253000, 854253900, 854254800,
    854255700, 854256600, 854257500, 854258400, 854259300, 854260200,
    854261100, 854262000, 854262900, 854263800, 854264700, 854265600,
    854266500, 854267400, 854268300, 854269200, 854270100, 854271000,
    854271900, 854272800, 854273700, 854274600, 854275500, 854276400,
    854277300, 854278200, 854279100, 854280000, 854280900, 854281800,
    854282700, 854283600, 854284500, 854285400, 854286300, 854287200,
    854288100, 854289000, 854289900, 854290800, 854291700, 854292600,
    854293500, 854294400, 854295300, 854296200, 854297100, 854298000,
    854298900, 854299800, 854328600, 854329500, 854330400, 854331300,
    854332200, 854333100, 854334000, 854334900, 854335800, 854336700,
    854337600, 854338500, 854339400, 854340300, 854341200, 854342100,
    854343000, 854343900, 854344800, 854345700, 854346600, 854347500,
    854348400, 854349300, 854350200, 854351100, 854352000, 854352900,
    854353800, 854354700, 854355600, 854356500, 854357400, 854358300,
    854359200, 854360100, 854361000, 854361900, 854362800, 854363700,
    854364600, 854365500, 854366400, 854367300, 854368200, 854369100,
    854370000, 854370900, 854371800, 854372700, 854373600, 854374500,
    854375400, 854376300, 854377200, 854378100, 854379000, 854379900,
    854380800, 854381700, 854382600, 854383500, 854384400, 854385300,
    854386200, 854387100, 854388000, 854388900, 854389800, 854390700,
    854391600, 854392500, 854393400, 854394300, 854395200, 854396100,
    854397000, 854397900, 854398800, 854399700, 854400600, 854401500,
    854402400, 854403300, 854404200, 854405100, 854406000, 854406900,
    854407800, 854408700, 854409600, 854410500, 854411400, 854412300,
    854413200, 854414100, 854415000, 854415900, 854416800, 854417700,
    854418600, 854419500, 854420400, 854421300, 854422200, 854423100,
    854424000, 854424900, 854425800, 854426700, 854427600, 854428500,
    854429400, 854430300, 854431200, 854432100, 854433000, 854433900,
    854434800, 854435700, 854436600, 854437500, 854438400, 854439300,
    854440200, 854441100, 854442000, 854442900, 854443800, 854444700,
    854445600, 854446500, 854447400, 854448300, 854449200, 854450100,
    854451000, 854451900, 854452800, 854453700, 854454600, 854455500,
    854456400, 854457300, 854458200, 854459100, 854460000, 854460900,
    854461800, 854462700, 854463600, 854464500, 854465400, 854466300,
    854467200, 854468100, 854469000, 854469900, 854470800, 854471700,
    854472600, 854473500, 854474400, 854475300, 854476200, 854477100,
    854478000, 854478900, 854479800, 854480700, 854481600, 854482500,
    854483400, 854484300, 854485200, 854486100, 854487000, 854487900,
    854488800, 854489700, 854490600, 854491500, 854492400, 854493300,
    854494200, 854495100, 854496000, 854496900, 854497800, 854498700,
    854499600, 854500500, 854501400, 854502300, 854503200, 854504100,
    854505000, 854505900, 854506800, 854507700, 854508600, 854509500,
    854510400, 854511300, 854512200, 854513100, 854514000, 854514900,
    854515800, 854516700, 854517600, 854518500, 854519400, 854520300,
    854521200, 854522100, 854523000, 854523900, 854524800, 854525700,
    854526600, 854527500, 854528400, 854529300, 854530200, 854531100,
    854532000, 854532900, 854533800, 854534700, 854535600, 854536500,
    854537400, 854538300, 854539200, 854540100, 854541000, 854541900,
    854542800, 854543700, 854544600, 854545500, 854546400, 854547300,
    854548200, 854549100, 854550000, 854550900, 854551800, 854552700,
    854553600, 854554500, 854555400, 854556300, 854557200, 854558100,
    854559000, 854559900, 854560800, 854561700, 854562600, 854563500,
    854564400, 854565300, 854566200, 854567100, 854568000, 854568900,
    854569800, 854570700, 854571600, 854572500, 854573400, 854574300,
    854575200, 854576100, 854577000, 854577900, 854578800, 854579700,
    854580600, 854581500, 854582400, 854583300, 854584200, 854585100,
    854586000, 854586900, 854587800, 854588700, 854589600, 854590500,
    854591400, 854592300, 854593200, 854594100, 854595000, 854595900,
    854596800, 854597700, 854598600, 854599500, 854600400, 854601300,
    854602200, 854603100, 854604000, 854604900, 854605800, 854606700,
    854607600, 854608500, 854609400, 854610300, 854611200, 854612100,
    854613000, 854613900, 854614800, 854615700, 854616600, 854617500,
    854618400, 854619300, 854620200, 854621100, 854622000, 854622900,
    854623800, 854624700, 854625600, 854626500, 854627400, 854628300,
    854629200, 854630100, 854631000, 854631900, 854632800, 854633700,
    854634600, 854635500, 854636400, 854637300, 854638200, 854639100,
    854640000, 854640900, 854641800, 854642700, 854643600, 854644500,
    854645400, 854646300, 854647200, 854648100, 854649000, 854649900,
    854650800, 854651700, 854652600, 854653500, 854654400, 854655300,
    854656200, 854657100, 854658000, 854658900, 854659800, 854660700,
    854661600, 854662500, 854663400, 854664300, 854665200, 854666100,
    854667000, 854667900, 854668800, 854669700, 854670600, 854671500,
    854672400, 854673300, 854674200, 854675100, 854676000, 854676900,
    854677800, 854678700, 854679600, 854680500, 854681400, 854682300,
    854683200, 854684100, 854685000, 854685900, 854686800, 854687700,
    854688600, 854689500, 854690400, 854691300, 854692200, 854693100,
    854694000, 854694900, 854695800, 854696700, 854697600, 854698500,
    854699400, 854700300, 854701200, 854702100, 854703000, 854703900,
    854704800, 854705700, 854706600, 854707500, 854708400, 854709300,
    854710200, 854711100, 854712000, 854712900, 854713800, 854714700,
    854715600, 854716500, 854717400, 854718300, 854719200, 854720100,
    854721000, 854721900, 854722800, 854723700, 854724600, 854725500,
    854726400, 854727300, 854728200, 854729100, 854730000, 854730900,
    854731800, 854732700, 854733600, 854734500, 854735400, 854736300,
    854737200, 854738100, 854739000, 854739900, 854740800, 854741700,
    854742600, 854743500, 854744400, 854745300, 854746200, 854747100,
    854748000, 854748900, 854749800, 854750700, 854751600, 854752500,
    854753400, 854754300, 854755200, 854756100, 854757000, 854757900,
    854758800, 854759700, 854760600, 854761500, 854762400, 854763300,
    854764200, 854765100, 854766000, 854766900, 854767800, 854768700,
    854769600, 854770500, 854771400, 854772300, 854773200, 854774100,
    854775000, 854775900, 854776800, 854777700, 854778600, 854779500,
    854780400, 854781300, 854782200, 854783100, 854784000, 854784900,
    854785800, 854786700, 854787600, 854788500, 854789400, 854790300,
    854791200, 854792100, 854793000, 854793900, 854794800, 854795700,
    854796600, 854797500, 854798400, 854799300, 854800200, 854801100,
    854802000, 854802900, 854803800, 854804700, 854805600, 854806500,
    854807400, 854808300, 854809200, 854810100, 854811000, 854811900,
    854812800, 854813700, 854814600, 854815500, 854816400, 854817300,
    854818200, 854819100, 854820000, 854820900, 854821800, 854822700,
    854823600, 854824500, 854825400, 854826300, 854827200, 854828100,
    854829000, 854829900, 854830800, 854831700, 854832600, 854833500,
    854834400, 854835300, 854836200, 854837100, 854838000, 854838900,
    854839800, 854840700, 854841600, 854842500, 854843400, 854844300,
    854845200, 854846100, 854847000, 854847900, 854848800, 854849700,
    854850600, 854851500, 854852400, 854853300, 854854200, 854855100,
    854856000, 854856900, 854857800, 854858700, 854859600, 854860500,
    854861400, 854862300, 854863200, 854864100, 854865000, 854865900,
    854866800, 854867700, 854868600, 854869500, 854870400, 854871300,
    854872200, 854873100, 854874000, 854874900, 854875800, 854876700,
    854877600, 854878500, 854879400, 854880300, 854881200, 854882100,
    854883000, 854883900, 854884800, 854885700, 854886600, 854887500,
    854888400, 854889300, 854890200, 854891100, 854892000, 854892900,
    854893800, 854894700, 854895600, 854896500, 854897400, 854898300,
    854899200, 854900100, 854901000, 854901900, 854902800, 854903700,
    854904600, 854905500, 854906400, 854907300, 854908200, 854909100,
    854910000, 854910900, 854911800, 854912700, 854913600, 854914500,
    854915400, 854916300, 854917200, 854918100, 854919000, 854919900,
    854920800, 854921700, 854922600, 854923500, 854924400, 854925300,
    854926200, 854927100, 854928000, 854928900, 854929800, 854930700,
    854931600, 854932500, 854933400, 854934300, 854935200, 854936100,
    854937000, 854937900, 854938800, 854939700, 854940600, 854941500,
    854942400, 854943300, 854944200, 854945100, 854946000, 854946900,
    854947800, 854948700, 854949600, 854950500, 854951400, 854952300,
    854953200, 854954100, 854955000, 854955900, 854956800, 854957700,
    854958600, 854959500, 854960400, 854961300, 854962200, 854963100,
    854964000, 854964900, 854965800, 854966700, 854967600, 854968500,
    854969400, 854970300, 854971200, 854972100, 854973000, 854973900,
    854974800, 854975700, 854976600, 854977500, 854978400, 854979300,
    854980200, 854981100, 854982000, 854982900, 854983800, 854984700,
    854985600, 854986500, 854987400, 854988300, 854989200, 854990100,
    854991000, 854991900, 854992800, 854993700, 854994600, 854995500,
    854996400, 854997300, 854998200, 854999100, 855000000, 855000900,
    855001800, 855002700, 855003600, 855004500, 855005400, 855006300,
    855007200, 855008100, 855009000, 855009900, 855010800, 855011700,
    855012600, 855013500, 855014400, 855015300, 855016200, 855017100,
    855018000, 855018900, 855019800, 855020700, 855021600, 855022500,
    855023400, 855024300, 855025200, 855026100, 855027000, 855027900,
    855028800, 855029700, 855030600, 855031500, 855032400, 855033300,
    855034200, 855035100, 855036000, 855036900, 855037800, 855038700,
    855039600, 855040500, 855041400, 855042300, 855043200, 855044100,
    855045000, 855045900, 855046800, 855047700, 855048600, 855049500,
    855050400, 855051300, 855052200, 855053100, 855054000, 855054900,
    855055800, 855056700, 855057600, 855058500, 855059400, 855060300,
    855061200, 855062100, 855063000, 855063900, 855064800, 855065700,
    855066600, 855067500, 855068400, 855069300, 855070200, 855071100,
    855072000, 855072900, 855073800, 855074700, 855075600, 855076500,
    855077400, 855078300, 855079200, 855080100, 855081000, 855081900,
    855082800, 855083700, 855084600, 855085500, 855086400, 855087300,
    855088200, 855089100, 855090000, 855090900, 855091800, 855092700,
    855093600, 855094500, 855095400, 855096300, 855097200, 855098100,
    855099000, 855099900, 855100800, 855101700, 855102600, 855103500,
    855104400, 855105300, 855106200, 855107100, 855108000, 855108900,
    855109800, 855110700, 855111600, 855112500, 855113400, 855114300,
    855115200, 855116100, 855117000, 855117900, 855118800, 855119700,
    855120600, 855121500, 855122400, 855123300, 855124200, 855125100,
    855126000, 855126900, 855127800, 855128700, 855129600, 855130500,
    855131400, 855132300, 855133200, 855134100, 855135000, 855135900,
    855136800, 855137700, 855138600, 855139500, 855140400, 855141300,
    855142200, 855143100, 855144000, 855144900, 855145800, 855146700,
    855147600, 855148500, 855149400, 855150300, 855151200, 855152100,
    855153000, 855153900, 855154800, 855155700, 855156600, 855157500,
    855158400, 855159300, 855160200, 855161100, 855162000, 855162900,
    855163800, 855164700, 855165600, 855166500, 855167400, 855168300,
    855169200, 855170100, 855171000, 855171900, 855172800, 855173700,
    855174600, 855175500, 855176400, 855177300, 855178200, 855179100,
    855180000, 855180900, 855181800, 855182700, 855183600, 855184500,
    855185400, 855186300, 855187200, 855188100, 855189000, 855189900,
    855190800, 855191700, 855192600, 855193500, 855194400, 855195300,
    855196200, 855197100, 855198000, 855198900, 855199800, 855200700,
    855201600, 855202500, 855203400, 855204300, 855205200, 855206100,
    855207000, 855207900, 855208800, 855209700, 855210600, 855211500,
    855212400, 855213300, 855214200, 855215100, 855216000, 855216900,
    855217800, 855218700, 855219600, 855220500, 855221400, 855222300,
    855223200, 855224100, 855225000, 855225900, 855226800, 855227700,
    855228600, 855229500, 855230400, 855231300, 855232200, 855233100,
    855234000, 855234900, 855235800, 855236700, 855237600, 855238500,
    855239400, 855240300, 855241200, 855242100, 855243000, 855243900,
    855244800, 855245700, 855246600, 855247500, 855248400, 855249300,
    855250200, 855251100, 855252000, 855252900, 855253800, 855254700,
    855255600, 855256500, 855257400, 855258300, 855259200, 855260100,
    855261000, 855261900, 855262800, 855263700, 855264600, 855265500,
    855266400, 855267300, 855268200, 855269100, 855270000, 855270900,
    855271800, 855272700, 855273600, 855274500, 855275400, 855276300,
    855277200, 855278100, 855279000, 855279900, 855280800, 855281700,
    855282600, 855283500, 855284400, 855285300, 855286200, 855287100,
    855288000, 855288900, 855289800, 855290700, 855291600, 855292500,
    855293400, 855294300, 855295200, 855296100, 855297000, 855297900,
    855298800, 855299700, 855300600, 855301500, 855302400, 855303300,
    855304200, 855305100, 855306000, 855306900, 855307800, 855308700,
    855309600, 855310500, 855311400, 855312300, 855313200, 855314100,
    855315000, 855315900, 855316800, 855317700, 855318600, 855319500,
    855320400, 855321300, 855322200, 855323100, 855324000, 855324900,
    855325800, 855326700, 855327600, 855328500, 855329400, 855330300,
    855331200, 855332100, 855333000, 855333900, 855334800, 855335700,
    855336600, 855337500, 855338400, 855339300, 855340200, 855341100,
    855342000, 855342900, 855343800, 855344700, 855345600, 855346500,
    855347400, 855348300, 855349200, 855350100, 855351000, 855351900,
    855352800, 855353700, 855354600, 855355500, 855356400, 855357300,
    855358200, 855359100, 855360000, 855360900, 855361800, 855362700,
    855363600, 855364500, 855365400, 855366300, 855367200, 855368100,
    855369000, 855369900, 855370800, 855371700, 855372600, 855373500,
    855374400, 855375300, 855376200, 855377100, 855378000, 855378900,
    855379800, 855380700, 855381600, 855382500, 855383400, 855384300,
    855385200, 855386100, 855387000, 855387900, 855388800, 855389700,
    855390600, 855391500, 855392400, 855393300, 855394200, 855395100,
    855396000, 855396900, 855397800, 855398700, 855399600, 855400500,
    855401400, 855402300, 855403200, 855404100, 855405000, 855405900,
    855406800, 855407700, 855408600, 855409500, 855410400, 855411300,
    855412200, 855413100, 855414000, 855414900, 855415800, 855416700,
    855417600, 855418500, 855419400, 855420300, 855421200, 855422100,
    855423000, 855423900, 855424800, 855425700, 855426600, 855427500,
    855428400, 855429300, 855430200, 855431100, 855432000, 855432900,
    855433800, 855434700, 855435600, 855436500, 855437400, 855438300,
    855439200, 855440100, 855441000, 855441900, 855442800, 855443700,
    855444600, 855445500, 855446400, 855447300, 855448200, 855449100,
    855450000, 855450900, 855451800, 855452700, 855453600, 855454500,
    855455400, 855456300, 855457200, 855458100, 855459000, 855459900,
    855460800, 855461700, 855462600, 855463500, 855464400, 855465300,
    855466200, 855467100, 855468000, 855468900, 855469800, 855470700,
    855471600, 855472500, 855473400, 855474300, 855475200, 855476100,
    855477000, 855477900, 855478800, 855479700, 855480600, 855481500,
    855482400, 855483300, 855484200, 855485100, 855486000, 855486900,
    855487800, 855488700, 855489600, 855490500, 855491400, 855492300,
    855493200, 855494100, 855495000, 855495900, 855496800, 855497700,
    855498600, 855499500, 855500400, 855501300, 855502200, 855503100,
    855504000, 855504900, 855505800, 855506700, 855507600, 855508500,
    855509400, 855510300, 855511200, 855512100, 855513000, 855513900,
    855514800, 855515700, 855516600, 855517500, 855518400, 855519300,
    855520200, 855521100, 855522000, 855522900, 855523800, 855524700,
    855525600, 855526500, 855527400, 855528300, 855529200, 855530100,
    855531000, 855531900, 855532800, 855533700, 855534600, 855535500,
    855536400, 855537300, 855538200, 855539100, 855540000, 855540900,
    855541800, 855542700, 855543600, 855544500, 855545400, 855546300,
    855547200, 855548100, 855549000, 855549900, 855550800, 855551700,
    855552600, 855553500, 855554400, 855555300, 855556200, 855557100,
    855558000, 855558900, 855559800, 855560700, 855561600, 855562500,
    855563400, 855564300, 855565200, 855566100, 855567000, 855567900,
    855568800, 855569700, 855570600, 855571500, 855572400, 855573300,
    855574200, 855575100, 855576000, 855576900, 855577800, 855578700,
    855579600, 855580500, 855581400, 855582300, 855583200, 855584100,
    855585000, 855585900, 855586800, 855587700, 855588600, 855589500,
    855590400, 855591300, 855592200, 855593100, 855594000, 855594900,
    855595800, 855596700, 855597600, 855598500, 855599400, 855600300,
    855601200, 855602100, 855603000, 855603900, 855604800, 855605700,
    855606600, 855607500, 855608400, 855609300, 855610200, 855611100,
    855612000, 855612900, 855613800, 855614700, 855615600, 855616500,
    855617400, 855618300, 855619200, 855620100, 855621000, 855621900,
    855622800, 855623700, 855624600, 855625500, 855626400, 855627300,
    855628200, 855629100, 855630000, 855630900, 855631800, 855632700,
    855633600, 855634500, 855635400, 855636300, 855637200, 855638100,
    855639000, 855639900, 855640800, 855641700, 855642600, 855643500,
    855644400, 855645300, 855646200, 855647100, 855648000, 855648900,
    855649800, 855650700, 855651600, 855652500, 855653400, 855654300,
    855655200, 855656100, 855657000, 855657900, 855658800, 855659700,
    855660600, 855661500, 855662400, 855663300, 855664200, 855665100,
    855666000, 855666900, 855667800, 855668700, 855669600, 855670500,
    855671400, 855672300, 855673200, 855674100, 855675000, 855675900,
    855676800, 855677700, 855678600, 855679500, 855680400, 855681300,
    855682200, 855683100, 855684000, 855684900, 855685800, 855686700,
    855687600, 855688500, 855689400, 855690300, 855691200, 855692100,
    855693000, 855693900, 855694800, 855695700, 855696600, 855697500,
    855698400, 855699300, 855700200, 855701100, 855702000, 855702900,
    855703800, 855704700, 855705600, 855706500, 855707400, 855708300,
    855709200, 855710100, 855711000, 855711900, 855712800, 855713700,
    855714600, 855715500, 855716400, 855717300, 855718200, 855719100,
    855720000, 855720900, 855721800, 855722700, 855723600, 855724500,
    855725400, 855726300, 855727200, 855728100, 855729000, 855729900,
    855730800, 855731700, 855732600, 855733500, 855734400, 855735300,
    855736200, 855737100, 855738000, 855738900, 855739800, 855740700,
    855741600, 855742500, 855743400, 855744300, 855745200, 855746100,
    855747000, 855747900, 855748800, 855749700, 855750600, 855751500,
    855752400, 855753300, 855754200, 855755100, 855756000, 855756900,
    855757800, 855758700, 855759600, 855760500, 855761400, 855762300,
    855763200, 855764100, 855765000, 855765900, 855766800, 855767700,
    855768600, 855769500, 855770400, 855771300, 855772200, 855773100,
    855774000, 855774900, 855775800, 855776700, 855777600, 855778500,
    855779400, 855780300, 855781200, 855782100, 855783000, 855783900,
    855784800, 855785700, 855786600, 855787500, 855788400, 855789300,
    855790200, 855791100, 855792000, 855792900, 855793800, 855794700,
    855795600, 855796500, 855797400, 855798300, 855799200, 855800100,
    855801000, 855801900, 855802800, 855803700, 855804600, 855805500,
    855806400, 855807300, 855808200, 855809100, 855810000, 855810900,
    855811800, 855812700, 855813600, 855814500, 855815400, 855816300,
    855817200, 855818100, 855819000, 855819900, 855820800, 855821700,
    855822600, 855823500, 855824400, 855825300, 855826200, 855827100,
    855828000, 855828900, 855829800, 855830700, 855831600, 855832500,
    855833400, 855834300, 855835200, 855836100, 855837000, 855837900,
    855838800, 855839700, 855840600, 855841500, 855842400, 855843300,
    855844200, 855845100, 855846000, 855846900, 855847800, 855848700,
    855849600, 855850500, 855851400, 855852300, 855853200, 855854100,
    855855000, 855855900, 855856800, 855857700, 855858600, 855859500,
    855860400, 855861300, 855862200, 855863100, 855864000, 855864900,
    855865800, 855866700, 855867600, 855868500, 855869400, 855870300,
    855871200, 855872100, 855873000, 855873900, 855874800, 855875700,
    855876600, 855877500, 855878400, 855879300, 855880200, 855881100,
    855882000, 855882900, 855883800, 855884700, 855885600, 855886500,
    855887400, 855888300, 855889200, 855890100, 855891000, 855891900,
    855892800, 855893700, 855894600, 855895500, 855896400, 855897300,
    855898200, 855899100, 855900000, 855900900, 855901800, 855902700,
    855903600, 855904500, 855905400, 855906300, 855907200, 855908100,
    855909000, 855909900, 855910800, 855911700, 855912600, 855913500,
    855914400, 855915300, 855916200, 855917100, 855918000, 855918900,
    855919800, 855920700, 855921600, 855922500, 855923400, 855924300,
    855925200, 855926100, 855927000, 855927900, 855928800, 855929700,
    855930600, 855931500, 855932400, 855933300, 855934200, 855935100,
    855936000, 855936900, 855937800, 855938700, 855939600, 855940500,
    855941400, 855942300, 855943200, 855944100, 855945000, 855945900,
    855946800, 855947700, 855948600, 855949500, 855950400, 855951300,
    855952200, 855953100, 855954000, 855954900, 855955800, 855956700,
    855957600, 855958500, 855959400, 855960300, 855961200, 855962100,
    855963000, 855963900, 855964800, 855965700, 855966600, 855967500,
    855968400, 855969300, 855970200, 855971100, 855972000, 855972900,
    855973800, 855974700, 855975600, 855976500, 855977400, 855978300,
    855979200, 855980100, 855981000, 855981900, 855982800, 855983700,
    855984600, 855985500, 855986400, 855987300, 855988200, 855989100,
    855990000, 855990900, 855991800, 855992700, 855993600, 855994500,
    855995400, 855996300, 855997200, 855998100, 855999000, 855999900,
    856000800, 856001700, 856002600, 856003500, 856004400, 856005300,
    856006200, 856007100, 856008000, 856008900, 856009800, 856010700,
    856011600, 856012500, 856013400, 856014300, 856015200, 856016100,
    856017000, 856017900, 856018800, 856019700, 856020600, 856021500,
    856022400, 856023300, 856024200, 856025100, 856026000, 856026900,
    856027800, 856028700, 856029600, 856030500, 856031400, 856032300,
    856033200, 856034100, 856035000, 856035900, 856036800, 856037700,
    856038600, 856039500, 856040400, 856041300, 856042200, 856043100,
    856044000, 856044900, 856045800, 856046700, 856047600, 856048500,
    856049400, 856050300, 856051200, 856052100, 856053000, 856053900,
    856054800, 856055700, 856056600, 856057500, 856058400, 856059300,
    856060200, 856061100, 856062000, 856062900, 856063800, 856064700,
    856065600, 856066500, 856067400, 856068300, 856069200, 856070100,
    856071000, 856071900, 856072800, 856073700, 856074600, 856075500,
    856076400, 856077300, 856078200, 856079100, 856080000, 856080900,
    856081800, 856082700, 856083600, 856084500, 856085400, 856086300,
    856087200, 856088100, 856089000, 856089900, 856090800, 856091700,
    856092600, 856093500, 856094400, 856095300, 856096200, 856097100,
    856098000, 856098900, 856099800, 856100700, 856101600, 856102500,
    856103400, 856104300, 856105200, 856106100, 856107000, 856107900,
    856108800, 856109700, 856110600, 856111500, 856112400, 856113300,
    856114200, 856115100, 856116000, 856116900, 856117800, 856118700,
    856119600, 856120500, 856121400, 856122300, 856123200, 856124100,
    856125000, 856125900, 856126800, 856127700, 856128600, 856129500,
    856130400, 856131300, 856132200, 856133100, 856134000, 856134900,
    856135800, 856136700, 856137600, 856138500, 856139400, 856140300,
    856141200, 856142100, 856143000, 856143900, 856144800, 856145700,
    856146600, 856147500, 856148400, 856149300, 856150200, 856151100,
    856152000, 856152900, 856153800, 856154700, 856155600, 856156500,
    856157400, 856158300, 856159200, 856160100, 856161000, 856161900,
    856162800, 856163700, 856164600, 856165500, 856166400, 856167300,
    856168200, 856169100, 856170000, 856170900, 856171800, 856172700,
    856173600, 856174500, 856175400, 856176300, 856177200, 856178100,
    856179000, 856179900, 856180800, 856181700, 856182600, 856183500,
    856184400, 856185300, 856186200, 856187100, 856188000, 856188900,
    856189800, 856190700, 856191600, 856192500, 856193400, 856194300,
    856195200, 856196100, 856197000, 856197900, 856198800, 856199700,
    856200600, 856201500, 856202400, 856203300, 856204200, 856205100,
    856206000, 856206900, 856207800, 856208700, 856209600, 856210500,
    856211400, 856212300, 856213200, 856214100, 856215000, 856215900,
    856216800, 856217700, 856218600, 856219500, 856220400, 856221300,
    856222200, 856223100, 856224000, 856224900, 856225800, 856226700,
    856227600, 856228500, 856229400, 856230300, 856231200, 856232100,
    856233000, 856233900, 856234800, 856235700, 856236600, 856237500,
    856238400, 856239300, 856240200, 856241100, 856242000, 856242900,
    856243800, 856244700, 856245600, 856246500, 856247400, 856248300,
    856249200, 856250100, 856251000, 856251900, 856252800, 856253700,
    856254600, 856255500, 856256400, 856257300, 856258200, 856259100,
    856260000, 856260900, 856261800, 856262700, 856263600, 856264500,
    856265400, 856266300, 856267200, 856268100, 856269000, 856269900,
    856270800, 856271700, 856272600, 856273500, 856274400, 856275300,
    856276200, 856277100, 856278000, 856278900, 856279800, 856280700,
    856281600, 856282500, 856283400, 856284300, 856285200, 856286100,
    856287000, 856287900, 856288800, 856289700, 856290600, 856291500,
    856292400, 856293300, 856294200, 856295100, 856296000, 856296900,
    856297800, 856298700, 856299600, 856300500, 856301400, 856302300,
    856303200, 856304100, 856305000, 856305900, 856306800, 856307700,
    856308600, 856309500, 856310400, 856311300, 856312200, 856313100,
    856314000, 856314900, 856315800, 856316700, 856317600, 856318500,
    856319400, 856320300, 856321200, 856322100, 856323000, 856323900,
    856324800, 856325700, 856326600, 856327500, 856328400, 856329300,
    856330200, 856331100, 856332000, 856332900, 856333800, 856334700,
    856335600, 856336500, 856337400, 856338300, 856339200, 856340100,
    856341000, 856341900, 856342800, 856343700, 856344600, 856345500,
    856346400, 856347300, 856348200, 856349100, 856350000, 856350900,
    856351800, 856352700, 856353600, 856354500, 856355400, 856356300,
    856357200, 856358100, 856359000, 856359900, 856360800, 856361700,
    856362600, 856363500, 856364400, 856365300, 856366200, 856367100,
    856368000, 856368900, 856369800, 856370700, 856371600, 856372500,
    856373400, 856374300, 856375200, 856376100, 856377000, 856377900,
    856378800, 856379700, 856380600, 856381500, 856382400, 856383300,
    856384200, 856385100, 856386000, 856386900, 856387800, 856388700,
    856389600, 856390500, 856391400, 856392300, 856393200, 856394100,
    856395000, 856395900, 856396800, 856397700, 856398600, 856399500,
    856400400, 856401300, 856402200, 856403100, 856404000, 856404900,
    856405800, 856406700, 856407600, 856408500, 856409400, 856410300,
    856411200, 856412100, 856413000, 856413900, 856414800, 856415700,
    856416600, 856417500, 856418400, 856419300, 856420200, 856421100,
    856422000, 856422900, 856423800, 856424700, 856425600, 856426500,
    856427400, 856428300, 856429200, 856430100, 856431000, 856431900,
    856432800, 856433700, 856434600, 856435500, 856436400, 856437300,
    856438200, 856439100, 856440000, 856440900, 856441800, 856442700,
    856443600, 856444500, 856445400, 856446300, 856447200, 856448100,
    856449000, 856449900, 856450800, 856451700, 856452600, 856453500,
    856454400, 856455300, 856456200, 856457100, 856458000, 856458900,
    856459800, 856460700, 856461600, 856462500, 856463400, 856464300,
    856465200, 856466100, 856467000, 856467900, 856468800, 856469700,
    856470600, 856471500, 856472400, 856473300, 856474200, 856475100,
    856476000, 856476900, 856477800, 856478700, 856479600, 856480500,
    856481400, 856482300, 856483200, 856484100, 856485000, 856485900,
    856486800, 856487700, 856488600, 856489500, 856490400, 856491300,
    856492200, 856493100, 856494000, 856494900, 856495800, 856496700,
    856497600, 856498500, 856499400, 856500300, 856501200, 856502100,
    856503000, 856503900, 856504800, 856505700, 856506600, 856507500,
    856508400, 856509300, 856510200, 856511100, 856512000, 856512900,
    856513800, 856514700, 856515600, 856516500, 856517400, 856518300,
    856519200, 856520100, 856521000, 856521900, 856522800, 856523700,
    856524600, 856525500, 856526400, 856527300, 856528200, 856529100,
    856530000, 856530900, 856531800, 856532700, 856533600, 856534500,
    856535400, 856536300, 856537200, 856538100, 856539000, 856539900,
    856540800, 856541700, 856542600, 856543500, 856544400, 856545300,
    856546200, 856547100, 856548000, 856548900, 856549800, 856550700,
    856551600, 856552500, 856553400, 856554300, 856555200, 856556100,
    856557000, 856557900, 856558800, 856559700, 856560600, 856561500,
    856562400, 856563300, 856564200, 856565100, 856566000, 856566900,
    856567800, 856568700, 856569600, 856570500, 856571400, 856572300,
    856573200, 856574100, 856575000, 856575900, 856576800, 856577700,
    856578600, 856579500, 856580400, 856581300, 856582200, 856583100,
    856584000, 856584900, 856585800, 856586700, 856587600, 856588500,
    856589400, 856590300, 856591200, 856592100, 856593000, 856593900,
    856594800, 856595700, 856596600, 856597500, 856598400, 856599300,
    856600200, 856601100, 856602000, 856602900, 856603800, 856604700,
    856605600, 856606500, 856607400, 856608300, 856609200, 856610100,
    856611000, 856611900, 856612800, 856613700, 856614600, 856615500,
    856616400, 856617300, 856618200, 856619100, 856620000, 856620900,
    856621800, 856622700, 856623600, 856624500, 856625400, 856626300,
    856627200, 856628100, 856629000, 856629900, 856630800, 856631700,
    856632600, 856633500, 856634400, 856635300, 856636200, 856637100,
    856638000, 856638900, 856639800, 856640700, 856641600, 856642500,
    856643400, 856644300, 856645200, 856646100, 856647000, 856647900,
    856648800, 856649700, 856650600, 856651500, 856652400, 856653300,
    856654200, 856655100, 856656000, 856656900, 856657800, 856658700,
    856659600, 856660500, 856661400, 856662300, 856663200, 856664100,
    856665000, 856665900, 856666800, 856667700, 856668600, 856669500,
    856670400, 856671300, 856672200, 856673100, 856674000, 856674900,
    856675800, 856676700, 856677600, 856678500, 856679400, 856680300,
    856681200, 856682100, 856683000, 856683900, 856684800, 856685700,
    856686600, 856687500, 856688400, 856689300, 856690200, 856691100,
    856692000, 856692900, 856693800, 856694700, 856695600, 856696500,
    856697400, 856698300, 856699200, 856700100, 856701000, 856701900,
    856702800, 856703700, 856704600, 856705500, 856706400, 856707300,
    856708200, 856709100, 856710000, 856710900, 856711800, 856712700,
    856713600, 856714500, 856715400, 856716300, 856717200, 856718100,
    856719000, 856719900, 856720800, 856721700, 856722600, 856723500,
    856724400, 856725300, 856726200, 856727100, 856728000, 856728900,
    856729800, 856730700, 856731600, 856732500, 856733400, 856734300,
    856735200, 856736100, 856737000, 856737900, 856738800, 856739700,
    856740600, 856741500, 856742400, 856743300, 856744200, 856745100,
    856746000, 856746900, 856747800, 856748700, 856749600, 856750500,
    856751400, 856752300, 856753200, 856754100, 856755000, 856755900,
    856756800, 856757700, 856758600, 856759500, 856760400, 856761300,
    856762200, 856763100, 856764000, 856764900, 856765800, 856766700,
    856767600, 856768500, 856769400, 856770300, 856771200, 856772100,
    856773000, 856773900, 856774800, 856775700, 856776600, 856777500,
    856778400, 856779300, 856780200, 856781100, 856782000, 856782900,
    856783800, 856784700, 856785600, 856786500, 856787400, 856788300,
    856789200, 856790100, 856791000, 856791900, 856792800, 856793700,
    856794600, 856795500, 856796400, 856797300, 856798200, 856799100,
    856800000, 856800900, 856801800, 856802700, 856803600, 856804500,
    856805400, 856806300, 856807200, 856808100, 856809000, 856809900,
    856810800, 856811700, 856812600, 856813500, 856814400, 856815300,
    856816200, 856817100, 856818000, 856818900, 856819800, 856820700,
    856821600, 856822500, 856823400, 856824300, 856825200, 856826100,
    856827000, 856827900, 856828800, 856829700, 856830600, 856831500,
    856832400, 856833300, 856834200, 856835100, 856836000, 856836900,
    856837800, 856838700, 856839600, 856840500, 856841400, 856842300,
    856843200, 856844100, 856845000, 856845900, 856846800, 856847700,
    856848600, 856849500, 856850400, 856851300, 856852200, 856853100,
    856854000, 856854900, 856855800, 856856700, 856857600, 856858500,
    856859400, 856860300, 856861200, 856862100, 856863000, 856863900,
    856864800, 856865700, 856866600, 856867500, 856868400, 856869300,
    856870200, 856871100, 856872000, 856872900, 856873800, 856874700,
    856875600, 856876500, 856877400, 856878300, 856879200, 856880100,
    856881000, 856881900, 856882800, 856883700, 856884600, 856885500,
    856886400, 856887300, 856888200, 856889100, 856890000, 856890900,
    856891800, 856892700, 856893600, 856894500, 856895400, 856896300,
    856897200, 856898100, 856899000, 856899900, 856900800, 856901700,
    856902600, 856903500, 856904400, 856905300, 856906200, 856907100,
    856908000, 856908900, 856909800, 856910700, 856911600, 856912500,
    856913400, 856914300, 856915200, 856916100, 856917000, 856917900,
    856918800, 856919700, 856920600, 856921500, 856922400, 856923300,
    856924200, 856925100, 856926000, 856926900, 856927800, 856928700,
    856929600, 856930500, 856931400, 856932300, 856933200, 856934100,
    856935000, 856935900, 856936800, 856937700, 856938600, 856939500,
    856940400, 856941300, 856942200, 856943100, 856944000, 856944900,
    856945800, 856946700, 856947600, 856948500, 856949400, 856950300,
    856951200, 856952100, 856953000, 856953900, 856954800, 856955700,
    856956600, 856957500, 856958400, 856959300, 856960200, 856961100,
    856962000, 856962900, 856963800, 856964700, 856965600, 856966500,
    856967400, 856968300, 856969200, 856970100, 856971000, 856971900,
    856972800, 856973700, 856974600, 856975500, 856976400, 856977300,
    856978200, 856979100, 856980000, 856980900, 856981800, 856982700,
    856983600, 856984500, 856985400, 856986300, 856987200, 856988100,
    856989000, 856989900, 856990800, 856991700, 856992600, 856993500,
    856994400, 856995300, 856996200, 856997100, 856998000, 856998900,
    856999800, 857000700, 857001600, 857002500, 857003400, 857004300,
    857005200, 857006100, 857007000, 857007900, 857008800, 857009700,
    857010600, 857011500, 857012400, 857013300, 857014200, 857015100,
    857016000, 857016900, 857017800, 857018700, 857019600, 857020500,
    857021400, 857022300, 857023200, 857024100, 857025000, 857025900,
    857026800, 857027700, 857028600, 857029500, 857030400, 857031300,
    857032200, 857033100, 857034000, 857034900, 857035800, 857036700,
    857037600, 857038500, 857039400, 857040300, 857041200, 857042100,
    857043000, 857043900, 857044800, 857045700, 857046600, 857047500,
    857048400, 857049300, 857050200, 857051100, 857052000, 857052900,
    857053800, 857054700, 857055600, 857056500, 857057400, 857058300,
    857059200, 857060100, 857061000, 857061900, 857062800, 857063700,
    857064600, 857065500, 857066400, 857067300, 857068200, 857069100,
    857070000, 857070900, 857071800, 857072700, 857073600, 857074500,
    857075400, 857076300, 857077200, 857078100, 857079000, 857079900,
    857080800, 857081700, 857082600, 857083500, 857084400, 857085300,
    857086200, 857087100, 857088000, 857088900, 857089800, 857090700,
    857091600, 857092500, 857093400, 857094300, 857095200, 857096100,
    857097000, 857097900, 857098800, 857099700, 857100600, 857101500,
    857102400, 857103300, 857104200, 857105100, 857106000, 857106900,
    857107800, 857108700, 857109600, 857110500, 857111400, 857112300,
    857113200, 857114100, 857115000, 857115900, 857116800, 857117700,
    857118600, 857119500, 857120400, 857121300, 857122200, 857123100,
    857124000, 857124900, 857125800, 857126700, 857127600, 857128500,
    857129400, 857130300, 857131200, 857132100, 857133000, 857133900,
    857134800, 857135700, 857136600, 857137500, 857138400, 857139300,
    857140200, 857141100, 857142000, 857142900, 857143800, 857144700,
    857145600, 857146500, 857147400, 857148300, 857149200, 857150100,
    857151000, 857151900, 857152800, 857153700, 857154600, 857155500,
    857156400, 857157300, 857158200, 857159100, 857160000, 857160900,
    857161800, 857162700, 857163600, 857164500, 857165400, 857166300,
    857167200, 857168100, 857169000, 857169900, 857170800, 857171700,
    857172600, 857173500, 904634100, 904635000, 904635900, 904636800,
    904637700, 904638600, 904639500, 904640400, 904641300, 904642200,
    904643100, 904644000, 904644900, 904645800, 904646700, 904647600,
    904648500, 904649400, 904650300, 904651200, 904652100, 904653000,
    904653900, 904654800, 904655700, 904656600, 904657500, 904658400,
    904659300, 904660200, 904661100, 904662000, 904662900, 904663800,
    904664700, 904665600, 904666500, 904667400, 904668300, 904669200,
    904670100, 904671000, 904671900, 904672800, 904673700, 904674600,
    904675500, 904676400, 904677300, 904678200, 904679100, 904680000,
    904680900, 904681800, 904682700, 904683600, 904684500, 904685400,
    904686300, 904687200, 904688100, 904689900, 904690800, 904691700,
    904692600, 904693500, 904694400, 904695300, 904696200, 904697100,
    904698000, 904698900, 904699800, 904700700, 904701600, 904702500,
    904703400, 904704300, 904705200, 904706100, 904707000, 904707900,
    904708800, 904709700, 904710600, 904711500, 904712400, 904713300,
    904714200, 904715100, 904716000, 904716900, 904717800, 904718700,
    904719600, 904720500, 904721400, 904722300, 904723200, 904724100,
    904725000, 904725900, 904726800, 904727700, 904728600, 904729500,
    904730400, 904731300, 904732200, 904733100, 904734000, 904734900,
    904735800, 904736700, 904737600, 904738500, 904739400, 904740300,
    904741200, 904742100, 904743000, 904743900, 904744800, 904745700,
    904746600, 904747500, 904748400, 904749300, 904750200, 904751100,
    904752000, 904752900, 904753800, 904754700, 904755600, 904756500,
    904757400, 904758300, 904759200, 904760100, 904761000, 904761900,
    904762800, 904763700, 904764600, 904765500, 904766400, 904767300,
    904768200, 904769100, 904770000, 904770900, 904771800, 904772700,
    904773600, 904774500, 904775400, 904776300, 904777200, 904778100,
    904779000, 904779900, 904780800, 904781700, 904782600, 904783500,
    904784400, 904785300, 904786200, 904787100, 904788000, 904788900,
    904789800, 904790700, 904791600, 904792500, 904793400, 904794300,
    904795200, 904796100, 904797000, 904797900, 904798800, 904799700,
    904800600, 904801500, 904802400, 904803300, 904804200, 904805100,
    904806000, 904806900, 904807800, 904808700, 904809600, 904810500,
    904811400, 904812300, 904813200, 904814100, 904815000, 904815900,
    904816800, 904817700, 904818600, 904819500, 904820400, 904821300,
    904822200, 904823100, 904824000, 904824900, 904825800, 904826700,
    904827600, 904828500, 904829400, 904830300, 904831200, 904832100,
    904833000, 904833900, 904834800, 904835700, 904836600, 904837500,
    904838400, 904839300, 904840200, 904841100, 904842000, 904842900,
    904843800, 904844700, 904845600, 904846500, 904847400, 904848300,
    904849200, 904850100, 904851000, 904851900, 904852800, 904853700,
    904854600, 904855500, 904856400, 904857300, 904858200, 904859100,
    904860000, 904860900, 904861800, 904862700, 904863600, 904864500,
    904865400, 904866300, 904867200, 904868100, 904869000, 904869900,
    904870800, 904871700, 904872600, 904873500, 904874400, 904875300,
    904876200, 904877100, 904878000, 904878900, 904879800, 904880700,
    904881600, 904882500, 904883400, 904884300, 904885200, 904886100,
    904887000, 904887900, 904888800, 904889700, 904890600, 904891500,
    904892400, 904893300, 904894200, 904895100, 904896000, 904896900,
    904897800, 904898700, 904899600, 904900500, 904901400, 904902300,
    904903200, 904904100, 904905000, 904905900, 904906800, 904907700,
    904908600, 904909500, 904910400, 904911300, 904912200, 904913100,
    904914000, 904914900, 904915800, 904916700, 904917600, 904918500,
    904919400, 904920300, 904921200, 904922100, 904923000, 904923900,
    904924800, 904925700, 904926600, 904927500, 904928400, 904929300,
    904930200, 904931100, 904932000, 904932900, 904933800, 904934700,
    904935600, 904936500, 904937400, 904938300, 904939200, 904940100,
    904941000, 904941900, 904942800, 904943700, 904944600, 904945500,
    904946400, 904947300, 904948200, 904949100, 904950000, 904950900,
    904951800, 904952700, 904953600, 904954500, 904955400, 904956300,
    904957200, 904958100, 904959000, 904959900, 904960800, 904961700,
    904962600, 904963500, 904964400, 904965300, 904966200, 904967100,
    904968000, 904968900, 904969800, 904970700, 904971600, 904972500,
    904973400, 904974300, 904975200, 904976100, 904977000, 904977900,
    904978800, 904979700, 904980600, 904981500, 904982400, 904983300,
    904984200, 904985100, 904986000, 904986900, 904987800, 904988700,
    904989600, 904990500, 904991400, 904992300, 904993200, 904994100,
    904995000, 904995900, 904996800, 904997700, 904998600, 904999500,
    905000400, 905001300, 905002200, 905003100, 905004000, 905004900,
    905005800, 905006700, 905007600, 905008500, 905009400, 905010300,
    905011200, 905012100, 905013000, 905013900, 905014800, 905015700,
    905016600, 905017500, 905018400, 905019300, 905020200, 905021100,
    905022000, 905022900, 905023800, 905024700, 905025600, 905026500,
    905027400, 905028300, 905029200, 905030100, 905031000, 905031900,
    905032800, 905033700, 905034600, 905035500, 905036400, 905037300,
    905038200, 905039100, 905040000, 905040900, 905041800, 905042700,
    905043600, 905044500, 905045400, 905046300, 905047200, 905048100,
    905049000, 905049900, 905050800, 905051700, 905052600, 905053500,
    905054400, 905055300, 905056200, 905057100, 905058000, 905058900,
    905059800, 905060700, 905061600, 905062500, 905063400, 905064300,
    905065200, 905066100, 905067000, 905067900, 905068800, 905069700,
    905070600, 905071500, 905072400, 905073300, 905074200, 905075100,
    905076000, 905076900, 905077800, 905078700, 905079600, 905080500,
    905081400, 905082300, 905083200, 905084100, 905085000, 905085900,
    905086800, 905087700, 905088600, 905089500, 905090400, 905091300,
    905092200, 905093100, 905094000, 905094900, 905095800, 905096700,
    905097600, 905098500, 905099400, 905100300, 905101200, 905102100,
    905103000, 905103900, 905104800, 905105700, 905106600, 905107500,
    905108400, 905109300, 905110200, 905111100, 905112000, 905112900,
    905113800, 905114700, 905115600, 905116500, 905117400, 905118300,
    905119200, 905120100, 905121000, 905121900, 905122800, 905123700,
    905124600, 905125500, 905126400, 905127300, 905128200, 905129100,
    905130000, 905130900, 905131800, 905132700, 905133600, 905134500,
    905135400, 905136300, 905137200, 905138100, 905139000, 905139900,
    905140800, 905141700, 905142600, 905143500, 905144400, 905145300,
    905146200, 905147100, 905148000, 905148900, 905149800, 905150700,
    905151600, 905152500, 905153400, 905154300, 905155200, 905156100,
    905157000, 905157900, 905158800, 905159700, 905160600, 905161500,
    905162400, 905163300, 905164200, 905165100, 905166000, 905166900,
    905167800, 905168700, 905169600, 905170500, 905171400, 905172300,
    905173200, 905174100, 905175000, 905175900, 905176800, 905177700,
    905178600, 905179500, 905180400, 905181300, 905182200, 905183100,
    905184000, 905184900, 905185800, 905186700, 905187600, 905188500,
    905189400, 905190300, 905191200, 905192100, 905193000, 905193900,
    905194800, 905195700, 905196600, 905197500, 905198400, 905199300,
    905200200, 905201100, 905202000, 905202900, 905203800, 905204700,
    905205600, 905206500, 905207400, 905208300, 905209200, 905210100,
    905211000, 905211900, 905212800, 905213700, 905214600, 905215500,
    905216400, 905217300, 905218200, 905219100, 905220000, 905220900,
    905221800, 905222700, 905223600, 905224500, 905225400, 905226300,
    905227200, 905228100, 905229000, 905229900, 905230800, 905231700,
    905232600, 905233500, 905234400, 905235300, 905236200, 905237100,
    905238000, 905238900, 905239800, 905240700, 905241600, 905242500,
    905243400, 905244300, 905245200, 905246100, 905247000, 905247900,
    905248800, 905249700, 905250600, 905251500, 905252400, 905253300,
    905254200, 905255100, 905256000, 905256900, 905257800, 905258700,
    905259600, 905260500, 905261400, 905262300, 905263200, 905264100,
    905265000, 905265900, 905266800, 905267700, 905268600, 905269500,
    905270400, 905271300, 905272200, 905273100, 905274000, 905274900,
    905275800, 905276700, 905277600, 905278500, 905279400, 905280300,
    905281200, 905282100, 905283000, 905283900, 905284800, 905285700,
    905286600, 905287500, 905288400, 905289300, 905290200, 905291100,
    905292000, 905292900, 905293800, 905294700, 905295600, 905296500,
    905297400, 905298300, 905299200, 905300100, 905301000, 905301900,
    905302800, 905303700, 905304600, 905305500, 905306400, 905307300,
    905308200, 905309100, 905310000, 905310900, 905311800, 905312700,
    905313600, 905314500, 905315400, 905316300, 905317200, 905318100,
    905319000, 905319900, 905320800, 905321700, 905322600, 905323500,
    905324400, 905325300, 905326200, 905327100, 905328000, 905328900,
    905329800, 905330700, 905331600, 905332500, 905333400, 905334300,
    905335200, 905336100, 905337000, 905337900, 905338800, 905339700,
    905340600, 905341500, 905342400, 905343300, 905344200, 905345100,
    905346000, 905346900, 905347800, 905348700, 905349600, 905350500,
    905351400, 905352300, 905353200, 905354100, 905355000, 905355900,
    905356800, 905357700, 905358600, 905359500, 905360400, 905361300,
    905362200, 905363100, 905364000, 905364900, 905365800, 905366700,
    905367600, 905368500, 905369400, 905370300, 905371200, 905372100,
    905373000, 905373900, 905374800, 905375700, 905376600, 905377500,
    905378400, 905379300, 905380200, 905381100, 905382000, 905382900,
    905383800, 905384700, 905385600, 905386500, 905387400, 905388300,
    905389200, 905390100, 905391000, 905391900, 905392800, 905393700,
    905394600, 905395500, 905396400, 905397300, 905398200, 905399100,
    905400000, 905400900, 905401800, 905402700, 905403600, 905404500,
    905405400, 905406300, 905407200, 905408100, 905409000, 905409900,
    905410800, 905411700, 905412600, 905413500, 905414400, 905415300,
    905416200, 905417100, 905418000, 905418900, 905419800, 905420700,
    905421600, 905422500, 905423400, 905424300, 905425200, 905426100,
    905427000, 905427900, 905428800, 905429700, 905430600, 905431500,
    905432400, 905433300, 905434200, 905435100, 905436000, 905436900,
    905437800, 905438700, 905439600, 905440500, 905441400, 905442300,
    905443200, 905444100, 905445000, 905445900, 905446800, 905447700,
    905448600, 905449500, 905450400, 905451300, 905452200, 905453100,
    905454000, 905454900, 905455800, 905456700, 905457600, 905458500,
    905459400, 905460300, 905461200, 905462100, 905463000, 905463900,
    905464800, 905465700, 905466600, 905467500, 905468400, 905469300,
    905470200, 905471100, 905472000, 905472900, 905473800, 905474700,
    905475600, 905476500, 905477400, 905478300, 905479200, 905480100,
    905481000, 905481900, 905482800, 905483700, 905484600, 905485500,
    905486400, 905487300, 905488200, 905489100, 905490000, 905490900,
    905491800, 905492700, 905493600, 905494500, 905495400, 905496300,
    905497200, 905498100, 905499000, 905499900, 905500800, 905501700,
    905502600, 905503500, 905504400, 905505300, 905506200, 905507100,
    905508000, 905508900, 905509800, 905510700, 905511600, 905512500,
    905513400, 905514300, 905515200, 905516100, 905517000, 905517900,
    905518800, 905519700, 905520600, 905521500, 905522400, 905523300,
    905524200, 905525100, 905526000, 905526900, 905527800, 905528700,
    905529600, 905530500, 905531400, 905532300, 905533200, 905534100,
    905535000, 905535900, 905536800, 905537700, 905538600, 905539500,
    905540400, 905541300, 905542200, 905543100, 905544000, 905544900,
    905545800, 905546700, 905547600, 905548500, 905549400, 905550300,
    905551200, 905552100, 905553000, 905553900, 905554800, 905555700,
    905556600, 905557500, 905558400, 905559300, 905560200, 905561100,
    905562000, 905562900, 905563800, 905564700, 905565600, 905566500,
    905567400, 905568300, 905569200, 905570100, 905571000, 905571900,
    905572800, 905573700, 905574600, 905575500, 905576400, 905577300,
    905578200, 905579100, 905580000, 905580900, 905581800, 905582700,
    905583600, 905584500, 905585400, 905586300, 905587200, 905588100,
    905589000, 905589900, 905590800, 905591700, 905592600, 905593500,
    905594400, 905595300, 905596200, 905597100, 905598000, 905598900,
    905599800, 905600700, 905601600, 905602500, 905603400, 905604300,
    905605200, 905606100, 905607000, 905607900, 905608800, 905609700,
    905610600, 905611500, 905612400, 905613300, 905614200, 905615100,
    905616000, 905616900, 905617800, 905618700, 905619600, 905620500,
    905621400, 905622300, 905623200, 905624100, 905625000, 905625900,
    905626800, 905627700, 905628600, 905629500, 905630400, 905631300,
    905632200, 905633100, 905634000, 905634900, 905635800, 905636700,
    905637600, 905638500, 905639400, 905640300, 905641200, 905642100,
    905643000, 905643900, 905644800, 905645700, 905646600, 905647500,
    905648400, 905649300, 905650200, 905651100, 905652000, 905652900,
    905653800, 905654700, 905655600, 905656500, 905657400, 905658300,
    905659200, 905660100, 905661000, 905661900, 905662800, 905663700,
    905664600, 905665500, 905666400, 905667300, 905668200, 905669100,
    905670000, 905670900, 905671800, 905672700, 905673600, 905674500,
    905675400, 905676300, 905677200, 905678100, 905679000, 905679900,
    905680800, 905681700, 905682600, 905683500, 905684400, 905685300,
    905686200, 905687100, 905688000, 905688900, 905689800, 905690700,
    905691600, 905692500, 905693400, 905694300, 905695200, 905696100,
    905697000, 905697900, 905698800, 905699700, 905700600, 905701500,
    905702400, 905703300, 905704200, 905705100, 905706000, 905706900,
    905707800, 905708700, 905709600, 905710500, 905711400, 905712300,
    905713200, 905714100, 905715000, 905715900, 905716800, 905717700,
    905718600, 905719500, 905720400, 905721300, 905722200, 905723100,
    905724000, 905724900, 905725800, 905726700, 905727600, 905728500,
    905729400, 905730300, 905731200, 905732100, 905733000, 905733900,
    905734800, 905735700, 905736600, 905737500, 905738400, 905739300,
    905740200, 905741100, 905742000, 905742900, 905743800, 905744700,
    905745600, 905746500, 905747400, 905748300, 905749200, 905750100,
    905751000, 905751900, 905752800, 905753700, 905754600, 905755500,
    905756400, 905757300, 905758200, 905759100, 905760000, 905760900,
    905761800, 905762700, 905763600, 905764500, 905765400, 905766300,
    905767200, 905768100, 905769000, 905769900, 905770800, 905771700,
    905772600, 905773500, 905774400, 905775300, 905776200, 905777100,
    905778000, 905778900, 905779800, 905780700, 905781600, 905782500,
    905783400, 905784300, 905785200, 905786100, 905787000, 905787900,
    905788800, 905789700, 905790600, 905791500, 905792400, 905793300,
    905794200, 905795100, 905796000, 905796900, 905797800, 905798700,
    905799600, 905800500, 905801400, 905802300, 905803200, 905804100,
    905805000, 905805900, 905806800, 905807700, 905808600, 905809500,
    905810400, 905811300, 905812200, 905813100, 905814000, 905814900,
    905815800, 905816700, 905817600, 905818500, 905819400, 905820300,
    905821200, 905822100, 905823000, 905823900, 905824800, 905825700,
    905826600, 905827500, 905828400, 905829300, 905830200, 905831100,
    905832000, 905832900, 905833800, 905834700, 905835600, 905836500,
    905837400, 905838300, 905839200, 905840100, 905841000, 905841900,
    905842800, 905843700, 905844600, 905845500, 905846400, 905847300,
    905848200, 905849100, 905850000, 905850900, 905851800, 905852700,
    905853600, 905854500, 905855400, 905856300, 905857200, 905858100,
    905859000, 905859900, 905860800, 905861700, 905862600, 905863500,
    905864400, 905865300, 905866200, 905867100, 905868000, 905868900,
    905869800, 905870700, 905871600, 905872500, 905873400, 905874300,
    905875200, 905876100, 905877000, 905877900, 905878800, 905879700,
    905880600, 905881500, 905882400, 905883300, 905884200, 905885100,
    905886000, 905886900, 905887800, 905888700, 905889600, 905890500,
    905891400, 905892300, 905893200, 905894100, 905895000, 905895900,
    905896800, 905897700, 905898600, 905899500, 905900400, 905901300,
    905902200, 905903100, 905904000, 905904900, 905905800, 905906700,
    905907600, 905908500, 905909400, 905910300, 905911200, 905912100,
    905913000, 905913900, 905914800, 905915700, 905916600, 905917500,
    905918400, 905919300, 905920200, 905921100, 905922000, 905922900,
    905923800, 905924700, 905925600, 905926500, 905927400, 905928300,
    905929200, 905930100, 905931000, 905931900, 905932800, 905933700,
    905934600, 905935500, 905936400, 905937300, 905938200, 905939100,
    905940000, 905940900, 905941800, 905942700, 905943600, 905944500,
    905945400, 905946300, 905947200, 905948100, 905949000, 905949900,
    905950800, 905951700, 905952600, 905953500, 905954400, 905955300,
    905956200, 905957100, 905958000, 905958900, 905959800, 905960700,
    905961600, 905962500, 905963400, 905964300, 905965200, 905966100,
    905967000, 905967900, 905968800, 905969700, 905970600, 905971500,
    905972400, 905973300, 905974200, 905975100, 905976000, 905976900,
    905977800, 905978700, 905979600, 905980500, 905981400, 905982300,
    905983200, 905984100, 905985000, 905985900, 905986800, 905987700,
    905988600, 905989500, 905990400, 905991300, 905992200, 905993100,
    905994000, 905994900, 905995800, 905996700, 905997600, 905998500,
    905999400, 906000300, 906001200, 906002100, 906003000, 906003900,
    906004800, 906005700, 906006600, 906007500, 906008400, 906009300,
    906010200, 906011100, 906012000, 906012900, 906013800, 906014700,
    906015600, 906016500, 906017400, 906018300, 906019200, 906020100,
    906021000, 906021900, 906022800, 906023700, 906024600, 906025500,
    906026400, 906027300, 906028200, 906029100, 906030000, 906030900,
    906031800, 906032700, 906033600, 906034500, 906035400, 906036300,
    906037200, 906038100, 906039000, 906039900, 906040800, 906041700,
    906042600, 906043500, 906044400, 906045300, 906046200, 906047100,
    906048000, 906048900, 906049800, 906050700, 906051600, 906052500,
    906053400, 906054300, 906055200, 906056100, 906057000, 906057900,
    906058800, 906059700, 906060600, 906061500, 906062400, 906063300,
    906064200, 906065100, 906066000, 906066900, 906067800, 906068700,
    906069600, 906070500, 906071400, 906072300, 906073200, 906074100,
    906075000, 906075900, 906076800, 906077700, 906078600, 906079500,
    906080400, 906081300, 906082200, 906083100, 906084000, 906084900,
    906085800, 906086700, 906087600, 906088500, 906089400, 906090300,
    906091200, 906092100, 906093000, 906093900, 906094800, 906095700,
    906096600, 906097500, 906098400, 906099300, 906100200, 906101100,
    906102000, 906102900, 906103800, 906104700, 906105600, 906106500,
    906107400, 906108300, 906109200, 906110100, 906111000, 906111900,
    906112800, 906113700, 906114600, 906115500, 906116400, 906117300,
    906118200, 906119100, 906120000, 906120900, 906121800, 906122700,
    906123600, 906124500, 906125400, 906126300, 906127200, 906128100,
    906129000, 906129900, 906130800, 906131700, 906132600, 906133500,
    906134400, 906135300, 906136200, 906137100, 906138000, 906138900,
    906139800, 906140700, 906141600, 906142500, 906143400, 906144300,
    906145200, 906146100, 906147000, 906147900, 906148800, 906149700,
    906150600, 906151500, 906152400, 906153300, 906154200, 906155100,
    906156000, 906156900, 906157800, 906158700, 906159600, 906160500,
    906161400, 906162300, 906163200, 906164100, 906165000, 906165900,
    906166800, 906167700, 906168600, 906169500, 906170400, 906171300,
    906172200, 906173100, 906174000, 906174900, 906175800, 906176700,
    906177600, 906178500, 906179400, 906180300, 906181200, 906182100,
    906183000, 906183900, 906184800, 906185700, 906186600, 906187500,
    906188400, 906189300, 906190200, 906191100, 906192000, 906192900,
    906193800, 906194700, 906195600, 906196500, 906197400, 906198300,
    906199200, 906200100, 906201000, 906201900, 906202800, 906203700,
    906204600, 906205500, 906206400, 906207300, 906208200, 906209100,
    906210000, 906210900, 906211800, 906212700, 906213600, 906214500,
    906215400, 906216300, 906217200, 906218100, 906219000, 906219900,
    906220800, 906221700, 906222600, 906223500, 906224400, 906225300,
    906226200, 906227100, 906228000, 906228900, 906229800, 906230700,
    906231600, 906232500, 906233400, 906234300, 906235200, 906236100,
    906237000, 906237900, 906238800, 906239700, 906240600, 906241500,
    906242400, 906243300, 906244200, 906245100, 906246000, 906246900,
    906247800, 906248700, 906249600, 906250500, 906251400, 906252300,
    906253200, 906254100, 906255000, 906255900, 906256800, 906257700,
    906258600, 906259500, 906260400, 906261300, 906262200, 906263100,
    906264000, 906264900, 906265800, 906266700, 906267600, 906268500,
    906269400, 906270300, 906271200, 906272100, 906273000, 906273900,
    906274800, 906275700, 906276600, 906277500, 906278400, 906279300,
    906280200, 906281100, 906282000, 906282900, 906283800, 906284700,
    906285600, 906286500, 906287400, 906288300, 906289200, 906290100,
    906291000, 906291900, 906292800, 906293700, 906294600, 906295500,
    906296400, 906297300, 906298200, 906299100, 906300000, 906300900,
    906301800, 906302700, 906303600, 906304500, 906305400, 906306300,
    906307200, 906308100, 906309000, 906309900, 906310800, 907373242,
    907374132, 907375034, 907375932, 907376837, 907377740, 907378638,
    907379539, 907380434, 907381340, 907382234, 907383135, 907384036,
    907384936, 907385834, 907386740, 907387634, 907388539, 907389435,
    907390335, 907391240, 907392136, 907393050, 907393941, 907394836,
    907395740, 907396641, 907397536, 907398436, 907399341, 907400237,
    907401136, 907402041, 907402941, 907403843, 907404736, 907405641,
    907406541, 907407436, 907408337, 907409237, 907410142, 907411036,
    907411936, 907412844, 907413742, 907414640, 907415536, 907416437,
    907417342, 907418237, 907419142, 907420038, 907420938, 907421837,
    907422737, 907423640, 907424542, 907425438, 907426341, 907427242,
    907428142, 907429042, 907429939, 907430838, 907431744, 907432642,
    907433544, 907434440, 907435339, 907436239, 907437138, 907438039,
    907438941, 907439839, 907440746, 907441639, 907442540, 907443447,
    907444342, 907445249, 907446146, 907447046, 907447941, 907448840,
    907449741, 907450641, 907451541, 907452446, 907453349, 907454249,
    907455148, 907456048, 907456942, 907457852, 907458754, 907459640,
    907460537, 907461435, 907462330, 907463231, 907464134, 907465033,
    907465938, 907466834, 907467735, 907468640, 907469535, 907470434,
    907471339, 907472236, 907473140, 907474035, 907474939, 907475835,
    907476735, 907477640, 907478535, 907479441, 907480341, 907481240,
    907482151, 907483042, 907483942, 907484836, 907485735, 907486635,
    907487536, 907488452, 907489336, 907490236, 907491136, 907492041,
    907492936, 907493836, 907494737, 907495666, 907496542, 907497438,
    907498336, 907499237, 907500142, 907501036, 907501936, 907502844,
    907503736, 907504638, 907505538, 907506444, 907507331, 907508231,
    907509131, 907510036, 907510936, 907511831, 907512735, 907513631,
    907514530, 907515436, 907516336, 907517231, 907518135, 907519032,
    907519935, 907520831, 907521736, 907522630, 907523536, 907524431,
    907525331, 907526231, 907527137, 907528037, 907528937, 907529836,
    907530737, 907531637, 907532531, 907533432, 907534336, 907535232,
    907536135, 907537030, 907537937, 907538836, 907539736, 907540631,
    907541534, 907542439, 907543334, 907544235, 907545134, 907546033,
    907546932, 907547832, 907548734, 907549632, 907550541, 907551434,
    907552337, 907553232, 907554138, 907555032, 907555932, 907556832,
    907557732, 907558633, 907559537, 907560432, 907561334, 907562232,
    907563132, 907564033, 907564938, 907565833, 907566732, 907567632,
    907568539, 907569432, 907570337, 907571232, 907572135, 907573033,
    907573932, 907574832, 907575732, 907576632, 907577537, 907578437,
    907579332, 907580234, 907581131, 907582032, 907582932, 907583838,
    907584731, 907585637, 907586531, 907587438, 907588331, 907589231,
    907590131, 907591031, 907591931, 907592832, 907593732, 907595550,
    907596433, 907597332, 907598240, 907599138, 907600032, 907600933,
    907601832, 907602737, 907603637, 907604533, 907605437, 907606337,
    907607232, 907608138, 907609037, 907609938, 907610832, 907611733,
    907612632, 907613532, 907614582, 907615332, 907616238, 907617132,
    907618032, 907618932, 907619832, 907620737, 907621632, 907622537,
    907623432, 907624333, 907625233, 907626134, 907627040, 907627932,
    907628837, 907629732, 907630637, 907631533, 907632436, 907633345,
    907634233, 907635131, 907636033, 907636933, 907637838, 907638732,
    907639633, 907640532, 907641437, 907642338, 907643232, 907644133,
    907645032, 907645934, 907646838, 907647732, 907648633, 907649533,
    907650432, 907651332, 907652238, 907653138, 907654038, 907654938,
    907655832, 907656738, 907657632, 907658532, 907659434, 907660332,
    907661246, 907662137, 907663036, 907663932, 907664834, 907665733,
    907666637, 907667537, 907668432, 907669332, 907670238, 907671132,
    907672037, 907672937, 907673832, 907674733, 907675632, 907676532,
    907677463, 907678332, 907679237, 907680132, 907681032, 907681933,
    907682832, 907683733, 907684632, 907685535, 907686438, 907687332,
    907688231, 907689131, 907690037, 907690932, 907691831, 907692736,
    907693633, 907694531, 907695437, 907696332, 907697237, 907698137,
    907699031, 907699931, 907700836, 907701731, 907702632, 907703531,
    907704431, 907705333, 907706236, 907707130, 907708030, 907708930,
    907709832, 907710738, 907711631, 907712532, 907713436, 907714332,
    907715232, 907716136, 907717031, 907717931, 907718835, 907719730,
    907720636, 907721530, 907722445, 907723339, 907724234, 907725133,
    907726037, 907726933, 907727838, 907728732, 907729637, 907730532,
    907731442, 907732333, 907733237, 907734137, 907735032, 907735933,
    907736834, 907737732, 907738634, 907739532, 907740432, 907741337,
    907742231, 907743132, 907744032, 907744931, 907745831, 907746736,
    907747644, 907748531, 907749437, 907750331, 907751236, 907752131,
    907753036, 907753931, 907754831, 907755736, 907756631, 907757536,
    907758436, 907759331, 907760231, 907761131, 907762035, 907762936,
    907763831, 907764730, 907765631, 907766535, 907767430, 907768330,
    907769230, 907770130, 907771030, 907771930, 907772835, 907773735,
    907774630, 907775530, 907776431, 907777335, 907778235, 907779135,
    907780030, 907780935, 907781830, 907782735, 907783634, 907784532,
    907785434, 907786329, 907787236, 907788130, 907789034, 907789930,
    907790829, 907791731, 907792634, 907793529, 907794430, 907795329,
    907796235, 907797130, 907798035, 907798930, 907799831, 907800735,
    907801631, 907802537, 907803436, 907804330, 907805229, 907806129,
    907807035, 907807929, 907808834, 907809734, 907810633, 907811546,
    907812438, 907813337, 907814232, 907815138, 907816038, 907816932,
    907817837, 907818733, 907819637, 907820537, 907821432, 907822332,
    907823234, 907824132, 907825031, 907825938, 907826837, 907827743,
    907828631, 907829533, 907830433, 907831333, 907832236, 907833131,
    907834067, 907834931, 907835832, 907836731, 907837636, 907838531,
    907839436, 907840346, 907841231, 907842131, 907843031, 907843931,
    907844831, 907845735, 907846636, 907847535, 907848435, 907849335,
    907850231, 907851130, 907852035, 907852938, 907853830, 907854730,
    907855632, 907856532, 907857433, 907858337, 907859237, 907860134,
    907861033, 907861937, 907862834, 907863737, 907864637, 907865536,
    907866431, 907867331, 907868233, 907869131, 907870037, 907870945,
    907871831, 907872736, 907873637, 907874533, 907875436, 907876336,
    907877232, 907878137, 907879031, 907879931, 907880831, 907881732,
    907882638, 907883539, 907884433, 907885332, 907886232, 907887136,
    907888032, 907888936, 907889833, 907890737, 911780267, 911781157,
    911782057, 911782957, 911783857, 911784757, 911785657, 911786557,
    911787457, 911788357, 911789257, 911790157, 911791057, 911791957,
    911792857, 911793757, 911794657, 911795557, 911796457, 911797357,
    911798257, 911799157, 911800057, 911800957, 911801857, 911802757,
    911803657, 911804557, 911805457, 911806357, 911807257, 911808157,
    911809057, 911809957, 911810857, 911811757, 911812657, 911813557,
    911814457, 911815357, 911816257, 911817157, 911818057, 911818957,
    911819857, 911820757, 911821657, 911822557, 911823457, 911824357,
    911825257, 911826157, 911827057, 911827957, 911828857, 911829757,
    911830657, 911831557, 911832457, 911833357, 911834257, 911835157,
    911836057, 911836957, 911837857, 911838757, 911839657, 911840557,
    911841457, 911842357, 911843257, 911844157, 911845057, 911845957,
    911846857, 911847757, 911848657, 911849555, 911850457, 911851357,
    911852257, 911853157, 911854057, 911854957, 911855860, 911856760,
    911857660, 911858557, 911859460, 911860360, 911861260, 911862160,
    911863060, 911863960, 911864860, 911865760, 911866667, 911867560,
    911868460, 911869360, 911870260, 911871160, 911872060, 911872960,
    911873860, 911874760, 911875660, 911876560, 911877461, 911878360,
    911879260, 911880160, 911881060, 911881960, 911882860, 911883760,
    911884660, 911885560, 911886460, 911887360, 911888260, 911889160,
    911890060, 911890960, 911891860, 911892760, 911893660, 911894560,
    911895460, 911896360, 911897260, 911898160, 911899062, 911899962,
    911900862, 911901762, 911902662, 911903562, 911904462, 911905362,
    911906262, 911907162, 911908062, 911908962, 911909862, 911910762,
    911911661, 911912562, 911913462, 911914362, 911915262, 911916162,
    911917062, 911917962, 911918862, 911919762, 911920662, 911921562,
    911922462, 911923362, 911924262, 911925162, 911926062, 911926962,
    911927862, 911928762, 911929662, 911930562, 911931462, 911932362,
    911933262, 911934162, 911935062, 911935962, 911936862, 911937762,
    911938662, 911939562, 911940462, 911941362, 911942262, 911943162,
    911944062, 911944962, 911945862, 911946762, 911947662, 911948562,
    911949462, 911950362, 911951262, 911952162, 911953067, 911953962,
    911954862, 911955762, 911956662, 911957562, 911958462, 911959362,
    911960262, 911961162, 911962062, 911962962, 911963862, 911964762,
    911965662, 911966562, 911967462, 911968362, 911969262, 911970162,
    911971062, 911971962, 911972862, 911973762, 911974662, 911975562,
    911976462, 911977362, 911978262, 911979162, 911980062, 911980962,
    911981862, 911982762, 911983662, 911984562, 911985462, 911986362,
    911987262, 911988162, 911989062, 911989962, 911990862, 911991762,
    911992662, 911993562, 911994462, 911995362, 911996262, 911997162,
    911998062, 911998962, 911999862, 912000762, 912001662, 912002562,
    912003462, 912004362, 912005262, 912006162, 912007062, 912007962,
    912008862, 912009762, 912010662, 912011562, 912012462, 912013362,
    912014262, 912015162, 912016062, 912016962, 912017862, 912018762,
    912019662, 912020562, 912021462, 912022362, 912023262, 912024162,
    912025062, 912025962, 912026862, 912027762, 912028662, 912029562,
    912030462, 912031362, 912032262, 912033162, 912034062, 912034962,
    912035862, 912036762, 912037662, 912038562, 912039472, 912040362,
    912041262, 912042162, 912043062, 912043962, 912044862, 912045762,
    912046662, 912047562, 912048462, 912049362, 912050262, 912051162,
    912052062, 912052962, 912053862, 912054762, 912055662, 912056562,
    912057462, 912058362, 912059262, 912060162, 912061062, 912061962,
    912062862, 912063762, 912064662, 912065562, 912066462, 912067362,
    912069128, 912070062, 912070962, 912071862, 912072762, 912073662,
    912074562, 912075462, 912076362, 912077262, 912078162, 912079062,
    912079962, 912080862, 912081762, 912082662, 912083562, 912084462,
    912085362, 912086262, 912087162, 912088062, 912088962, 912089862,
    912090762, 912091662, 912092562, 912093462, 912094362, 912095262,
    912096162, 912097062, 912097962, 912098862, 912099762, 912100662,
    912101562, 912102462, 912103362, 912104262, 912105162, 912106062,
    912106962, 912107862, 912108762, 912109662, 912110562, 912111462,
    912112362, 912113262, 912114162, 912115062, 912115962, 912116862,
    912117762, 912118662, 912119562, 912120462, 912121362, 912122262,
    912123162, 912124062, 912124962, 912125872, 912126762, 912127662,
    912128562, 912129462, 912130362, 912131262, 912132162, 912133062,
    912133962, 912134862, 912135762, 912136662, 912137562, 912138462,
    912139362, 912140262, 912141162, 912142062, 912142962, 912143862,
    912144762, 912145662, 912146562, 912147462, 912148362, 912149262,
    912150162, 912151062, 912151962, 912152862, 912153762, 912154662,
    912155562, 912156462, 912157362, 912158262, 912159162, 912160062,
    912160962, 912161862, 912162762, 912163662, 912164562, 912165462,
    912166362, 912167262, 912168162, 912169062, 912169962, 912170862,
    912171762, 912172662, 912173562, 912174462, 912175362, 912176262,
    912177162, 912178062, 912178962, 912179862, 912180762, 912181662,
    912182562, 912183462, 912184362, 912185262, 912186162, 912187062,
    912187962, 912188862, 912189762, 912190662, 912191562, 912192462,
    912193362, 912194262, 912195162, 912196062, 912196962, 912197862,
    912198762, 912199662, 912200562, 912201462, 912202362, 912203262,
    912204162, 912205062, 912205962, 912206862, 912207762, 912208662,
    912209562, 912210462, 912211362, 912212272, 912213162, 912214062,
    912214962, 912215862, 912216762, 912217662, 912218562, 912219462,
    912220362, 912221262, 912222162, 912223062, 912223962, 912224862,
    912225762, 912226662, 912227562, 912228462, 912229362, 912230262,
    912231162, 912232062, 912232962, 912233862, 912234762, 912235662,
    912236562, 912237462, 912238362, 912239262, 912240162, 912241062,
    912241962, 912242862, 912243762, 912244662, 912245562, 912246462,
    912247362, 912248262, 912249162, 912250062, 912250962, 912251862,
    912252762, 912253662, 912254562, 912255462, 912256362, 912257262,
    912258162, 912259062, 912259962, 912260862, 912261762, 912262662,
    912263562, 912264462, 912265362, 912266262, 912267162, 912268062,
    912268962, 912269862, 912270762, 912271662, 912272562, 912273462,
    912274362, 912275262, 912276162, 912277062, 912277962, 912278862,
    912279762, 912280662, 912281562, 912282462, 912283362, 912284262,
    912285162, 912286062, 912286962, 912287862, 912288762, 912289662,
    912290562, 912291462, 912292362, 912293262, 912294162, 912295062,
    912295962, 912296862, 912297762, 912298672, 912299562, 912300462,
    912301362, 912302262, 912303162, 912304062, 912304962, 912305862,
    912306762, 912307662, 912308562, 912309462, 912310362, 912311262,
    912312162, 912313062, 912313962, 912314862, 912315762, 912316662,
    912317562, 912318462, 912319356, 912320262, 912321162, 912322062,
    912322962, 912323862, 912324762, 912325662, 912326562, 912327462,
    938757947, 938813564, 938972137, 939003957, 939037502, 939185102,
    939228605, 939458142, 940206915, 940207822, 940209622, 940210522,
    940211422, 940212322, 940213222, 940214122, 940215022, 940216822,
    940218622, 940219522, 940220417, 940221322, 940223122, 940224020,
    940225795, 940226722, 940228522, 940229422, 940230322, 940231222,
    940232122, 940233922, 940234822, 940235722, 940236622, 940237522,
    940238422, 940239322, 940240222, 940246515, 940249222, 940257375,
    940258272, 940259170, 940260069, 940260976, 940261874, 940262774,
    940263669, 940264571, 940270862, 940271770, 940279817, 940283422,
    940286122, 940287022, 940287922, 940288822, 940289722, 940290622,
    940291522, 940420222, 940422022, 940424722, 940440922, 940445422,
    940449922, 940450822, 940452622, 940453522, 940454422, 940456222,
    940457122, 940458022, 940458922, 940459822, 940460722, 940461622,
    940462522, 940463422, 940464322, 940724547, 940725437, 940726337,
    940727237, 940728137, 940729037, 940729937, 940730837, 940731737,
    940732637, 940733537, 940734437, 940735337, 940736237, 940737137,
    940738037, 940738937, 940739837, 940740737, 940741637, 940742537,
    940743437, 940744337, 940745237, 940746137, 940747037, 940747937,
    940748837, 940749737, 940750637, 940751537, 940752437, 940753337,
    940755103, 940756037, 940756937, 940757837, 940758737, 940759637,
    940760537, 940761439, 940762337, 940763237, 940764137, 940765037,
    940765937, 940766837, 940767737, 940768637, 940769537, 940770437,
    940771337, 940772237, 940773137, 940774037, 940774937, 940775837,
    940776737, 940777637, 940778537, 940779437, 940780337, 940781237,
    940782137, 940783037, 940783937, 940784837, 940785737, 940786637,
    940787537, 940788437, 940789337, 940790237, 940791137, 940792037,
    940792937, 940793837, 940794737, 940795637, 940796537, 940797437,
    940798337, 940799237, 940800137, 940801037, 940801937, 940802837,
    940803737, 940804637, 940805537, 940806437, 940807337, 940808237,
    940809137, 940810037 ;
}
